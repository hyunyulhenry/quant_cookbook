"","SPY","IEV","EWJ","EEM","TLT","IEF","IYR","RWX","GLD","DBC"
"1",0.00212235483819123,-0.0056814470354658,0.0105634486272226,-0.0138089777070859,0.00606314442295375,0.0036283859050168,-0.000238122535192176,-0.00743650039460242,-0.01011555892928,-0.0260503050587256
"2",-0.00797616615140428,-0.0147621811294277,-0.0257840791300752,-0.0292382644144845,-0.00435264944621672,-0.00325455305176137,-0.0155039691262139,-0.0124342563723361,-0.0240065523436642,-0.0034512995305368
"3",0.00462505785007039,0.00164362834500564,0.00572253572691861,0.00725719012180659,0.00179373416960282,0.000725519952708087,-0.000242241519382569,-0.00338989013623814,0.00515210254785115,0.00519471605092869
"4",-0.000850250439833444,-0.00376383560049154,0.00640105341404884,-0.0223361655072509,0,-0.000241625017845748,0.0117532527075166,0.00161970411012868,0.00611769179894184,-0.00861317890472024
"5",0.00333185383113022,-0.00561872122315621,-0.0148410172356069,-0.00230329759424897,-0.00447651902474167,-0.00169178390223657,0.0159285448715216,-0.00565978108129528,-0.00427276924479103,-0.0147698688123383
"6",0.00438052067814776,0.0108136598205906,-0.00502142829521812,0.0126501433345514,-0.0058437181116715,-0.00266249523578876,0.0114341377918188,0.00325267589994183,0.000660191450734482,-0.00132265790941177
"7",0.00759715402776329,0.00905914380438233,0.012977654262998,0.0203336969156163,-0.00463587085246731,-0.00206404320428055,0.0034964852693331,0.00664608132280797,0.0253999171136414,0.0233996224013486
"8",-0.00195491429036387,0,0.00355853205057222,0.00357477449165522,0.00215850610712831,0.00194658047481866,0.0114984966606249,0.00257678539125261,-0.0032169375331168,-0.0228645994088241
"9",0.000419724192354476,-0.00057304824329707,0,-0.00418516439316152,-0.00306095299356002,-0.00194279866087899,0.00298501418550279,0.00706676333734224,0.0108116506243077,0.00883002834000157
"10",-0.00335622895000676,-0.00305809478065688,-0.000709148162663986,-0.0105519514238314,0.00307035119423937,0.00133831468790868,-0.00343391209739841,-0.00111624593135951,-0.00606642729991103,-0.0105032427762808
"11",0.00196451504111472,0.0107364911411358,0.00709716327695142,0.0179850132533814,-0.00272077042811147,-0.00157944223357942,0.00884477898830749,0.00973961024955017,0.0118856733660673,0.0150376039605462
"12",-0.00308078921929666,-0.00701852575518147,0,-0.00115424583911428,0.00238713446468308,0.00182486505287649,-0.0030739481740939,0.010278311948732,-0.00444442857142857,0.000871366900456527
"13",0.00294981649084236,0.00897792590611513,0.00563793367584275,0.0227532330831659,-0.00657572382122174,-0.00291462947491106,0.00285562622078328,0.00751315203843106,0.0240752866059424,0.0317805604448693
"14",0.0080529171210304,0.00511179600558109,0.0133145799163663,0.00869061932587689,-0.000114658458510775,0.000121826427972316,0.0136672140256091,0.00093170740976789,0.00155688923134556,-0.00843882505047222
"15",-0.0117400336575767,-0.0154451339250472,-0.0165973490401511,-0.0307572789044992,-0.0071903440947424,-0.0038963443820238,0.00595553165547646,-0.00589736158688503,-0.00419717070737846,-0.00893599478055107
"16",-0.000913958638936618,0.00277388619729968,0.000702927752839422,0.00613326450503893,-0.000805364687838428,-0.000122219315075833,0.0030155400881029,-0.00624540061248458,0.00171714023469072,0.0124515654514379
"17",-0.000562426957088857,0.00228937836540988,0.00351375549550559,-0.0132524430965038,-0.0021863081160356,-0.000733096116484866,0.0028947788506779,0.00612728098557302,-0.00623341144564171,-0.020356203459988
"18",0.00520975627008013,0.00532981302560187,0.00630267383024541,0.0154896664835846,0.0011528328306738,0.000977817344071097,0.00344267786464925,0.00405963517940289,0.00705662537243201,0.027705554222162
"19",0.00672290827199484,0.00511194143821414,-0.00417532450434566,0.00775909297911315,0.00840861183908359,0.00366709545627208,0.0113973095258864,0,0.00949861399099006,0.0105308029970261
"20",0.0059823412622575,0.00781788600721289,0.0132773618769466,0.0122480189860927,-0.00120484225647355,-0.000721096020748213,-0.000547218060078514,0.0113530302068443,0.00601571784619104,-0.00375161049023653
"21",0.00138306869815663,-0.000934605986404935,-0.00620689907498195,-0.00302503939292709,0.00126380958987471,0.00085621049210749,0.00711564741572834,0.0110720456488449,-0.0144127872675132,0.0129706315284444
"22",0.00027662460690081,-0.00327423655290127,-0.00763353448627713,0.000953849250799887,0.00137619303573433,0.00110057044765388,-0.000652021466787889,0.00304141699126781,0.000466692602157481,-0.00330437818714768
"23",0.000275724481370698,0.00656976193527181,0.00839171797977034,0.00987340000263726,0.00549633884997935,0.00280811068639153,0.0137043107551313,0.0103109727542583,0.00746389387230284,-0.00497302215289619
"24",0.00220865333901199,0.00372976539313519,-0.000693643549549372,-0.00385930099273324,0.00296097988774546,0.00219191605356484,0.0147000162874038,0.00405240375739147,-0.00246957860056218,-0.0120781760068096
"25",-0.00130846714880994,-0.0023223791723983,-0.0124914998459981,-0.00533792453258242,0.000795620028676725,0.000242973858452844,-0.0076136374241178,-0.000597976059040772,0.0137706953630217,0.0231870629732278
"26",-0.00744739017206775,-0.00595931686280271,0.0028111715201582,-0.0119449851553155,-0.00567345686755338,-0.00303661408258227,-0.0141714867859879,0.000598333848357502,0.00915760115190478,0.00618051849681645
"27",-0.00340426288464779,-0.00327819738511537,-0.000700785356489764,-0.00683301014310367,-0.00228202005450462,-0.00134072380076111,-0.0167532352453277,-0.00822062978989824,-0.00680588293379225,-0.0188371198035659
"28",0.0084350669567792,0.00977352256735409,0.0210378336471537,0.0158771923118854,-0.00217382087942752,-0.000731142424647779,0.0178076726966532,0.00813813313396716,0.00258867070469515,0.0183639546801622
"29",0.00656692990097851,0.012843145344263,0.016483502561536,0.0215332804796007,0.00951470076980976,0.00573835815185642,-0.00615586447707006,0.0165947142645049,0.00804992454738307,-0.0135245569450847
"30",0.00130515226998562,-0.00202127542937802,0.00810796746504328,0.000594920337946947,0.00295169350475621,0.00157704362551025,0.00825917372171392,0.00294110331554465,0.00060269697441484,0
"31",-0.000480291222614504,-0.000276345719207538,-0.000670091816536211,0.00229403426731922,0.00350979725290546,0.00109123331822802,-0.00344898850326691,-0.000733535898917448,-0.000752943788408844,0.0174491644849777
"32",0.00212708402943163,0.00349958807310791,-0.00335342141618133,0.00262722434384988,0.00225615442415505,0.0012104344485524,0.00843614648619351,0.00190797364020545,-0.015822829779644,-0.0110249158425911
"33",-0.000411141561985295,-0.00734191770007731,0.000672961455531862,0.00295815791524867,-0.00168805077046219,-0.00012165075553372,-0.00525534929064886,0.00322176900980553,0.0312356463400902,0.0214698305811687
"34",-0.0007529484591422,0.00286603530410812,0.00268993301217724,-0.0025284473772873,-0.00541229114787023,-0.0025385976482114,-0.00506716136696406,0.00627740276346822,-0.00296950268654794,0.013742936552138
"35",-0.00390764099820973,0.0025814158309363,0.00871910017145616,-0.00718192335541168,0.00714185002365864,0.00400132323481239,-0.0141961685093741,0.00681837709850708,0.00848844352975586,0.00637963267720099
"36",-0.000894484639078708,0.00505723257650148,0.006648870663025,-0.00042540488468068,0.0066418642666024,0.0031397055302802,-0.00648532507035171,-0.0080690587744835,0.00561129643220171,0.00277337747782158
"37",-0.039057911818374,-0.0539797589651595,-0.0237779997195946,-0.0813112101773937,0.0126352632133897,0.00842651461120059,-0.0324193345321695,-0.0368969497153717,-0.0395006472687415,-0.0189648488774585
"38",0.0102508936623875,0.0135396929246925,-0.00135329040260435,0.0250231500191431,-0.00452751185589384,-0.00346185874464677,0.00777632981289145,-0.00558096570895805,0.0163583387030521,0.0153039919303792
"39",-0.00298044613228909,-0.0131677865761087,-0.00474243921543993,-0.0143761011824965,-0.000634435668741107,0.000900894068910585,-0.00624087652201688,-0.0121339656036809,-0.00992784251228152,-0.00713994426755238
"40",-0.0130948820407214,-0.0130538223423906,-0.0163377949158395,-0.00926534596875328,0.00501341806506161,0.00324312229900436,-0.0206669177650952,-0.0188854332533552,-0.0320571406867212,-0.00918906513063011
"41",-0.00951882491150391,-0.0202802726485757,-0.0145329208160516,-0.0256479890148159,0.00166298720374014,0.000597341541918928,-0.0354435766774029,-0.0228480055468765,-0.0122429604809757,-0.0149191936410714
"42",0.0171094706175756,0.0276002791959264,0.0238765807448114,0.0439036793773289,-0.00298825015865445,-0.00131565120643606,0.0344494808358784,0.0281869443628027,0.0193866518353727,0.00941465989397505
"43",-0.00100237615288468,0.00194630887603853,-0.00205771841604041,-0.00609923213466057,0.00388554470673297,0.00179702612116039,-0.0142555778344917,0.011837814595115,0.00233828519600054,0.0137874316339257
"44",0.00845538929719192,0.0103921203866397,0.00893474676034223,0.0258288264705291,-0.000884899827255259,-0.000120070862838939,0.0160032050613381,0.00369457705078591,0.00279937778540984,0.00160000109706515
"45",0.000283990768656039,0.00288392299807483,0.000681296107118534,0.00178612247356358,-0.0105146047859809,-0.00561997114714918,0.012249821958167,0.0111964386500916,-0.00356704387870443,-0.0131789655455684
"46",0.00149181569209622,0.00383404043896163,0.00816876254923216,0.00490160926474981,0.00391542041851456,0.00276612277499222,0.00507162051216903,0.00712896540787922,0.00186775097276271,-0.00930789262729326
"47",-0.0194339529848233,-0.0244437308822566,-0.0182309316812997,-0.0290906946734778,0.00601651899175182,0.00443633819452205,-0.0263755260480876,-0.0191265782965131,-0.0100979022791097,-0.00776139923920816
"48",0.00744983664821675,0.00371937922979915,-0.00894089108085183,0.0082213996463949,-0.00454111880105834,-0.00131262165100066,0.0047110076735084,-0.0196531785542494,0.00345257370601737,0.00205841743606472
"49",0.00136439381968034,0.00477789241622006,0.00069412502489552,0.00815439476960855,-0.000110831483971618,-0.00107625314710302,0.0075027029776662,0.0117464222989827,0.000625602136778314,-0.00616274323701982
"50",-0.00280008131724463,0.0034937961555106,-0.000693643549549372,-0.00853801249608155,-0.000223536054364204,-0.000118665589326383,-0.00558492430364621,-0.00346377056960701,0.0100031728665209,0.00248040983341546
"51",0.0120551585124433,0.0149904973330299,0.0111033767470741,0.0219365530068458,-0.00211393182528685,-0.00131770693696465,0.0100629781599539,0.019485362266233,0.001856932751922,0.00494845688755019
"52",0.00549221494728402,0.00981403388292557,0.00892248211239877,0.00656378045720207,0.000556830922243901,0.00143828184344663,0.00324405784971127,0.0151373669027863,0.00818657733044725,0.00123089067396864
"53",0.0164574723223323,0.0245329850795801,0.0108843511171168,0.0299607704452685,0.00044696090071894,0.00143594885735299,0.0140869945467306,0.0227443743523146,0.00842658227791837,0.00163947728165459
"54",-0.000767661528157215,-0.00653891912286053,0.00134584084009148,-0.00427785120718527,-0.00791108943622765,-0.00334559843673443,-0.000796645258032691,-0.005890841857491,-0.000911546642357819,0.0163664913648924
"55",0.00146671460743408,0.00519146589935993,0.00134417541811938,0.00464005703573256,-0.00280873124696213,-0.0015592032839632,-0.000264015525573758,-0.000444381951905104,-0.00927615543564009,0.000402619932218462
"56",-0.00132504928910149,0.000737451822004243,-0.00536936136791577,-0.000598567991106691,0.00123896139924518,0.000841163234452269,-0.0155086352399035,-0.00340913928964537,0.0105908515551543,0.00442656260043939
"57",-0.00237463867980348,-0.00608222956638382,-0.00404840025328812,-0.00445030411881486,-0.00168581148953029,-0.000240637664685628,-0.00828443445884086,-0.00654353313353384,-0.00212635189102994,0.0028045321486756
"58",-0.00727942710823926,-0.00917954572881796,-0.00745252251999162,-0.0178804558497069,-0.00202868716150573,-0.000119778138517823,-0.0116483331355891,-0.00748539376289814,0.00532733662073093,0.00958850037405323
"59",0.00105718017456846,0.0103874095163914,0.00136504946009786,0.0198690166944311,-0.00135457649947812,-0.00144059304737743,0.00535730242056287,0.00829590944429404,-0.00605603303303415,0.0193905524746216
"60",0.000211718632761926,0.00342710258784806,-0.00681656670538833,-0.000171371992107483,-0.00192236462168849,-0.00120198560120965,0.00935391852372125,0.0127151568603869,0.00137084535046927,-0.0147516879941152
"61",0.00112655752060342,0.00359983160951161,-0.00549089021858618,0.00686667714845512,0.001659346252886,0.00111153115243345,0.0118494758302177,0.0053173865982763,0.00167325834113963,-0.00985019969883938
"62",0.0107627694881034,0.0129679101795244,0.00828170462817934,0.0163682063322272,-0.00124745219332456,-0.000844482930251189,0.00869564823080005,0.00573033717697014,-0.000303659842176507,-0.00397922538928086
"63",0.001113443862236,0.00254208637838649,0.00752926702828605,0.0062908471932468,0.00102167809181597,0.00157004690136153,-0.00655162737371817,-0.000876864017575585,0.0148867684980474,0.0111865837697289
"64",0.00271123234945692,0.00443776074955826,-0.00271750944657612,0.000917149464970235,-0.00374600806641179,-0.00253203455118234,0.000809212294691219,0.00438665850657571,0.000748435885299825,0.00197546276217331
"65",0.00138617182207845,-0.000991871460438332,-0.00136242605965198,0.00574623482636394,-0.00660979371922221,-0.0045954257951657,-0.000693221024568258,0.000145397400631797,-0.00493571634855339,-0.0102523310478511
"66",0.00117713128033348,0.00722028807430797,0.00341077438500492,0.00471954668250496,0.00298289641383898,0.00206566619030979,0.00254493762358221,0.00611380727748201,0.00946948759160504,0.0139442326305543
"67",-0.00408002471630187,-0.00394250357155157,-0.00407892131244625,-0.0092301576480246,-0.000686640496837421,-0.00121195937910901,-0.0133856816902801,-0.0111395064363944,-0.00119121493798613,-0.00157179448515576
"68",0.0044439343533007,0.00710665171022273,-0.00136502864824439,0.0167192972759918,0.0002284978180076,0.000970416612544156,-0.00526254103672041,0.00555920380988129,-0.00134174116452757,0.00590315003881492
"69",0.00456234891534102,0.00741413958928616,-0.00820251320691545,0.00490890979360059,-0.00308916397099235,-0.0016972528478173,0.0109348328047025,-0.00334632357876852,0.0126884314879365,0.00547739648670853
"70",0.00949633066192068,0.0117039976117963,0.0144728881349361,0.0118861717016479,0.00550996060435249,0.00109319220805304,-0.000233196151525839,0.0157660895113374,0.00825480591125038,-0.00778202330855171
"71",0.0026584270646075,0.00131475184029761,-0.00611404931401727,-0.00539078088836098,0.00559351008616105,0.00424602518622685,0.0143094491119062,-0.0054610486234753,-0.00584798228514671,-0.0101961268708496
"72",0.001223989762559,-0.000525043946775883,0.00136689449839378,-0.00744194304197887,0.00499481362343701,0.00229519098098518,-0.00355608061115087,-0.00173420445178063,0.00558819117647058,0.000396154335922549
"73",-0.000271479003905006,0,-0.00477813097111568,-0.00806830304201334,-0.00169472867200715,-0.000120956897947222,-0.00863222467036395,-0.00376335741437994,-0.0124305065412623,-0.00277227922738532
"74",0.00944059251763285,0.00796903061946175,0.0041152068025827,0.0119132133174236,-0.00260227574803484,-0.0010849723170977,0.0109137123585235,0.00624803398599094,0.0173256036920717,0.0138999306258629
"75",-0.00376816008539105,-0.00564732072804763,-0.0109288753716594,-0.00397851200956556,0.00363078457006338,0.00205170200451765,0.0084990958832476,-0.00216653407895862,-0.00640458543251454,0.00665883749617335
"76",0.000405411915245457,0.000174717471578711,-0.00138139130624471,-0.000162971292866132,0.00372981469503419,0.00192642848073765,-0.00683322144061282,-0.00723566970473943,-0.0077644152427655,-0.0136186866940441
"77",0.00918195706434632,0.0105704404061056,0.00553257619194913,0.0123928979787151,-0.00349030647210846,-0.000600204792663206,0.0013760510225338,0.009183482683911,0.00236226181770594,0.019723922310988
"78",0.00113723208839156,-0.00311165505497513,-0.00481430015824069,-0.00265772136689901,-0.00723325288526178,-0.00288676370634544,0.00137377067317779,-0.00548908767649403,-0.0150242453236743,-0.00696329557888986
"79",-0.00080233961460241,0.000259700014310527,-0.00552858371672771,-0.00500646041669217,-0.000227249309140087,0,-0.00331563102838583,-0.000725931996690576,0.0103184532532472,0.00506419748851039
"80",-0.00829226325219012,-0.0039009217342838,-0.00764446072803826,-0.0193147833762282,0.0104746204461088,0.00434217030591988,-0.0191602235813995,-0.00218015713070319,-0.00695680896852591,-0.00891469419041446
"81",0.00256260130802843,0.000261036847139851,0,0.00397206159562646,0.000723949793850265,0.0000483453927115907,-0.00526361182449586,-0.0033504255748662,-0.0059620513317663,0.00195550177609105
"82",0.00585165037666546,0.00539449858300833,0.00560246451473922,0.0198646892151604,-0.000564970669825748,-0.001205854482627,0.00823072858795704,0.020169812817457,-0.000449812552112516,-0.00780644828912236
"83",0.00541660994283544,-0.000865322462401452,0.00139270147481896,0.00840553494981022,-0.00226161785203183,-0.00108556277744509,0.00396575613143346,0.00286508748173842,0.0124511543683676,0.00472082218868608
"84",0.0037913401744456,0.012126497658171,0.00347718702147004,-0.00032058179557215,0.00407969472151115,0.00253721653728523,-0.00499545992092465,0.00628561591895083,0.0103719665245805,-0.00195784038455937
"85",0.00019889482245028,0,0.00485082990224139,0.00649425440611129,0.00270916300145951,0.000842886143124222,0.000934056229760172,0.00525289938824969,0.000879865057050289,-0.00470760579377849
"86",-0.00132541921592622,-0.00898608348890595,-0.00206892430402872,-0.0129840919289171,-0.00225214355345016,0,-0.00653217306927312,-0.012145451044643,-0.00542128937728936,-0.00630683405612698
"87",0.00271997312622929,0.00276386397667649,0.0124395346054402,0.0161406542820308,-0.00394798688084919,-0.00325088919923922,0.0116240972665291,0.00114387307203434,-0.00633470858874685,-0.00515664530307158
"88",-0.0104525564637009,-0.0201518831413005,-0.0150169384552497,-0.0244616730670175,0.00237895544663336,0.00253742999173867,-0.00998146399634059,-0.00756813279733126,-0.0214973619643007,-0.00398732915969924
"89",0.00855757066009888,0.01687440920081,0.00762286853376204,0.0254005686869998,-0.00350351246512159,-0.00204922103359684,0.0111372451955012,0.0141009845427646,0.00681813636363637,0.0148119473263204
"90",-0.00218776084110039,-0.00216048906061439,-0.00275106760484156,-0.00992458799659701,-0.00260827133474384,-0.00144871277598602,-0.0104350144637323,-0.0039733630213602,-0.00255828453987728,-0.00355029840873888
"91",0.000265998784142019,0.00259834422849736,-0.00827582337901067,0.00120306029185691,-0.000341147891411708,-0.000120575961113256,-0.0134738615084017,0.00284930094311009,0.00392278219557607,0.00989703519012286
"92",0.00684090644458224,0.00216006846614691,0.0020861892376951,0.0144975472101769,-0.000681676147225474,-0.000604141993891472,-0.00926383299678413,-0.00724417448258075,-0.0141268858712521,-0.00980004381165411
"93",-0.00197894091741069,-0.00172436592431247,-0.00832759603573918,-0.0036321094714088,-0.00409706099737794,-0.00266270829921611,-0.0179812362671461,-0.00887150180728025,-0.00823170756803993,0.00831350277362031
"94",0.00872406522999247,0.0125218186465905,-0.00279919708628318,0.00515096712373531,-0.0066277082764713,-0.00291219173792412,-0.00866686472246514,-0.00389735931653135,0.00707038140394678,-0.00157051832110122
"95",-0.000524113319638086,-0.00759071203903516,0,0.00181347295366008,0.0029912138880126,0.0013389760590643,0.0068955733608056,-0.00130439452177322,0.00228939265671824,0.00983104263365253
"96",-0.000786684964893758,0.00120299786015798,0.00982478733076642,0.000157131367967578,-0.00516121890538024,-0.0027949081359554,0.0103954175332859,0.000580020753876642,-0.00715701255236845,-0.014408109306017
"97",0.000131183118199374,0.00472108868529797,0.00138971318578474,-0.00157380044134237,-0.00288258831656696,-0.00195013547681444,-0.00786782014408194,0.00203076727295914,0.00521478551601784,0.00474108523167938
"98",-0.00905265797371546,-0.0105935130299306,-0.00485764798255295,-0.0240348196359494,0.000925518558194005,0.0013431644529609,-0.015249403913039,-0.0123025689089276,-0.0120537227333885,-0.00550522883832627
"99",0.00417088005447264,0.00682151114313778,-0.00418431437043032,0.0153415728567659,-0.00231041871975302,-0.00109713465233641,0.00631793761052424,0.000292741392376117,0.00293439382239402,0.0122577335130811
"100",0.00362569596282225,0.000428523135259873,0.0105045062029749,-0.00341990802406034,-0.000116330010013099,-0.0020756656586306,0.0305309304347514,-0.000585776757517142,0.00200181700025182,-0.0218748918446232
"101",0.00814464005283178,0.00488654191842497,0.00207879127072053,0.0102140010549032,0.00208437566438158,0.000978697908132764,0.0255641170973198,0.0063031044024453,-0.00537880743814345,0.00958467109811956
"102",-0.00104229356825192,0.00153572926680678,0.00968176585477165,0.00284362258960669,-0.00184835669194094,-0.000366233870316646,-0.00267895546288532,0.0180627390127408,0.012669962721416,0.00909802267606286
"103",0.00495712687915906,0.00894358011399699,0.00547960824917082,0.0249687085141439,-0.00525416838681347,-0.00430838526073551,-0.000466764758367044,0.00300418548259174,0.0137320870654245,0.00744810721222477
"104",0.000129701967523932,0.00303946401832511,0.00340587822522154,-0.00445687779336734,0.00455779326136319,0.001602492632514,0.00630955224479068,0.00699020539232831,0.00150510230267598,0.00894950605841682
"105",-0.00395876961403108,-0.00547107483769249,-0.00135755316700314,-0.00347406071131062,-0.00628131354031214,-0.0032008424542348,-0.0173016481861565,-0.00878288449343601,-0.00255482412752006,-0.00385662185426483
"106",-0.0107499364608572,-0.019803797772653,-0.00407892131244625,-0.0251740576099074,-0.00046782802741685,0.000494424824317052,-0.00626211530850163,-0.0195798392521699,0.00060269697441484,-0.00038718847866448
"107",-0.0180452300273917,-0.0231391551176165,-0.00409543974624027,-0.0154153122701323,-0.0179155491236713,-0.00999618049667372,-0.0309158934038625,-0.0236152857290732,-0.0173166982492577,0.00503486046064849
"108",0.0130112759089636,0.0142301890291019,0.0047976128104803,0.017674317317683,-0.000834945646363106,0.00186979880455085,0.016441376563695,0.00104533654531536,-0.0159362698150086,-0.0177263688049796
"109",0.00172190479734358,0.000435819810067795,-0.00136418080851974,0.00856453686221914,-0.00286354063629035,-0.00261268864661146,-0.0147263986292466,-0.00372854960385582,0.00747424466717161,0.0192232805596453
"110",-0.010905653325215,-0.0164634976537413,-0.0129782438596471,-0.0173769193330072,-0.014481754923155,-0.00711053878096701,-0.021073168154395,-0.0176643358064833,-0.00927355529861917,-0.00269446454548161
"111",0.0149682511328839,0.0172704617003778,0.00276803372271828,0.0200049487879173,0.011901364442205,0.00326614514971357,0.021526806160441,0.0118863659458568,0.00670828414066427,0.0127363633446651
"112",0.00638581078045908,0.00948964812643371,0.00138045945190224,0.0156895346495765,-0.0025202449215862,0.000250413379926373,-0.010291868468673,0.00135523093129097,0.00108475129528518,0.00952748724430674
"113",0.00569034057539231,0.0125055414391109,0.00895937692259241,0.0227855180651497,0.00685751218917763,0.00438236358517585,0.0151028812423089,0.00811273732363138,0.00386996916006099,0.00604001949708444
"114",-0.00117605079762051,0.00212927936610474,-0.00204928518371184,0.00090597809933346,-0.00203131209732332,-0.000498843490800094,-0.0148781778885561,-0.0033089662536856,0.00154200467361609,0
"115",0.00248534475428741,0.00144504543524793,-0.000684560398927059,0.00113201455145151,0.00933973639103636,0.00486366918534875,0.000990430859105773,0.00739462463042484,0.00816021592733862,-0.00975602421892541
"116",-0.0138972074365992,-0.012985987630718,-0.00684916573980365,-0.00851659384496517,-0.00806690896527396,-0.0032264896844395,-0.0178085385425711,-0.0112356796452635,-0.011759376370218,0.00113671378480618
"117",0.00555771395519877,0.0061054674010339,0.00482756013323149,0.0124661661078524,-0.00478378087627718,-0.00124542776769776,-0.00402958556532185,0.0037877848859651,-0.00231804979629191,-0.00454197639049791
"118",-0.00940914785959113,-0.00965825249949781,-0.00960858704466394,-0.0132132299356579,0.00648902840891918,0.00299226536816399,-0.00379260290766714,-0.00981142913405342,0.00340769837074673,-0.00228145187285711
"119",-0.00478214402757837,-0.00276163075156577,-0.00554407726304174,-0.00760804924166769,0.00549191411545147,0.00323234728467225,-0.0227155555255361,-0.0213412028090774,-0.00540288677682743,-0.0038110602241177
"120",-0.0102788794662315,-0.00519260263987698,0.00139365074198361,-0.00873978827196031,0.000237133941101142,0.000247881756367585,-0.00142831781103581,0.0023361390514125,-0.0125717988514669,-0.0114765510385546
"121",0.0142295236528327,0.0091346154839278,0.00208772590429351,0.0142307172884031,0.000949498580795405,-0.000124200711083655,0.0217165855627646,0.00310852039697851,0.000785900672522821,-0.00154803023238326
"122",-0.000133359998416904,0.00206890135442728,-0.00208337638544531,0.000228593610482442,-0.00023619756246307,-0.000619576494245266,-0.00390650861344022,0.00898493432604774,0.00926659366315663,-0.00310073611494466
"123",0.000332795991880852,0.00593606613352371,0.00974250871296767,0.00350701921699881,0.0103194378611846,0.00520627001206053,-0.00128968432229315,-0.002303023168716,0.000155539988934361,-0.00077756390523942
"124",0.00904073316747134,0.0116309102547412,0.0179185857439246,0.0202841044573383,0.00525673336178389,0.00152338709980682,0.0251870093395239,0.0110805620515233,0.011669519760519,0.00622568534584866
"125",0.00362344308847096,0.006086572153992,-0.00203116583233764,0.00796731172658705,-0.00609711685513614,-0.00296662235967871,-0.00466147952519047,0.000456350664309602,-0.0043063520904193,0.00116001076655725
"126",-0.00105086121150177,-0.0034452067399634,-0.00271359525328907,0.00443229934836298,-0.0112062667266896,-0.00557951501999843,0.0160754678604174,-0.00654208636489773,-0.00494284846904058,0.00926999570093279
"127",0.00525743253981603,0.00758880000932982,-0.00476171305520023,0.0171359987729978,-0.00405621925963473,-0.00236843018854194,-0.00211741641624075,0.0124045476708141,0.00838250569334065,0.00841948881502264
"128",0.000784421630519061,0.00343098009555143,0,0.00968909069923241,0.00359399591145482,0.00362368651411926,0.00374529307151694,-0.00862216206784183,0.00646548655273227,-0.0022770415146578
"129",-0.0142391313071289,-0.0146774173466412,0.0020503521677413,-0.0196935724158199,0.0169487992309301,0.00684875077099156,-0.0304726134564307,-0.0122063638930779,0.00351795672306299,0.00722704709078603
"130",0.00709009606728661,0.0131183803760544,-0.00341067039671283,0.00825466619980375,-0.010329068372637,-0.00346284343531322,0,0.00447975618613494,-0.00259105315361896,0.00226594368689348
"131",0.0157900274888354,0.0167086179038469,0.00684479010469952,0.0219534257246066,-0.00343886243221814,-0.00285387297406547,0.0125721733094175,0.00830360723608958,0.00886300400785434,0.0026375300692274
"132",0.00297946359515544,-0.00246509932357197,0.00475866207782749,0.0124070368972877,0.00273726123117823,0.00223979039753441,0.00950157809432994,0.00732068391602492,0.000151499552476508,0.00150315505542631
"133",-0.000128511625293481,-0.0023063048085098,-0.00202995623270441,-0.0098040566504235,0.00961302550461363,0.00397340425168768,-0.00552165360093892,-0.00408798599999149,-0.0031803574614625,-0.017636035275769
"134",-0.000516976216264009,-0.00132118349987298,-0.0054237383571436,-0.000777680718001883,-0.0021160374141449,-0.00210272563841019,-0.00643611305797975,-0.00881726018594953,-0.00106350653296861,-0.00611145817995895
"135",-0.00180937381787272,-0.00727507946593542,-0.00477170061118615,-0.0122442719389997,0.00376885562471463,0.00359455592459312,-0.00546152095165808,-0.00153346888472328,0.0132319847908744,0.011529517868204
"136",0.0038841747127456,0.0044135382650714,0.00479457890628354,0.00995971854253641,-0.000234686500699133,-0.000124135486219146,0.00331992092593048,0.00153582402307495,0.00585408259438247,0.00341949609782533
"137",-0.010124479053817,-0.0092029340989308,-0.00408994002323293,-0.00688182371236534,0.00903914904068959,0.00494133475372038,-0.0160378585017827,0.00076687033196543,0.00850619285162812,-0.000378725846339356
"138",0.00306187642854838,0.00317971831607222,0.00616022970577257,0.0289329062825907,-0.0016287999520429,-0.000368864429694304,-0.0174649319041688,-0.00766267605227922,-0.00162771525221317,-0.00454541746867632
"139",-0.017341227514907,-0.0212712345598042,-0.00340132731618448,-0.0342291772159689,0.00372876041800407,0.00270513645879977,-0.0256747274408309,-0.02007743830718,0,-0.00761027412690252
"140",0.00204929349029115,-0.00196052603185892,0.000682524730049039,0.00575114056106818,0.00197347871594844,0.00134866641025133,0.00135128165313758,0.00315211606127286,-0.00844818425302818,0.00881890096296867
"141",-0.0236794726561109,-0.0379159863285692,-0.0177352448100691,-0.0509649046240505,0.00834196467451087,0.00795988140597403,-0.0229420615387287,-0.0416340773961934,-0.0186846033278145,-0.0106421866674594
"142",-0.0196592566051441,-0.015178338242352,-0.00972227491988931,-0.012954847405439,0.00287203572081807,0.00194389802073847,-0.0276241919148704,-0.0186882172084319,-0.00365571961444877,0.00960418518193684
"143",0.0156429984519819,0.0208198641982129,0.0168302797463482,0.0327355927746129,-0.00286381075403497,-0.00254581516507946,0.0134945079848121,0.00818588839345802,0.00550363825080957,-0.0114154519572044
"144",-0.0112634536617956,0.00573948648774314,-0.004827412943186,-0.020466846675945,0.00723996539937577,0.00413331462211985,-0.0133148308930099,0.012261496108908,0.000304150842518558,0.00808306373567436
"145",0.00487244608969739,-0.000527132112596362,-0.00762318547098906,-0.00392212131784686,-0.00216570420217377,-0.00277189991288807,0.0156253192496554,-0.00965787185317302,0.002127967743913,-0.00152730162096215
"146",0.00799030191507666,0.00368897704491089,-0.00488834823728235,0.0110559869759697,0.00252501292727514,0.000731426619463793,0.0146849066229675,0.00495867252200277,-0.00060671924768696,0.0015296378393137
"147",-0.0257454081510448,-0.0175022068901207,-0.0140349519857694,-0.0431427138823994,0.00663994099534171,0.00645484286955256,-0.0368018071352125,-0.0149668306889765,0.0121414935823569,-0.0110728958450327
"148",0.0167597862349242,0.0115792673467332,0.0149465811135809,0.017847181292771,-0.00727807782749379,-0.00399330463813652,0.0260440300218061,0.001001506632335,-0.00254918270957627,-0.0138994995789665
"149",0.0106695401140731,0.00255351676402493,-0.00210398007030288,0.00746009474834608,-0.000801808240292856,-0.000120873423004708,0.00404474726443205,0.0158468515912125,-0.000601232739081525,0.00548151681725861
"150",0.013940518180924,0.0209028414607042,0.00843317174251856,0.0335876178754384,-0.0121543061878446,-0.0069261508018601,0.0362551896332204,0.0279144810328746,0.00436212375020517,-0.00155763343848836
"151",-0.0296337066985093,-0.0351858314956044,-0.0160280140095544,-0.0413586703520218,0.0013936773113854,0.00562742380826031,-0.00174291235585899,-0.0190095625426939,-0.0196195605640062,-0.00780031722738583
"152",-0.00467710761743922,-0.0141774257510432,-0.0141643410606317,-0.0173346848678908,-0.00231751905361288,-0.00145939582425436,-0.0331675435270334,-0.00749059575681787,0.0169569357921926,0.00353769611988386
"153",0.00359329272151876,-0.00018105272980895,0.00143681150591668,0.00987884217664403,0.00290386472565918,0.00158377324717729,-0.00416682671629309,-0.00459418223798436,-0.00465672224725844,-0.00705053381947773
"154",-0.0152861603065689,-0.00986059503186076,-0.00286932510624893,-0.0258521117636407,0.00266392659322934,0.00365042598823884,-0.0376564769915637,-0.0214272434283239,0.000452746741540944,0.0031557362828909
"155",-0.0137751033376641,-0.0244859612151852,-0.0165468193363462,-0.0392895442146558,-0.00358056020805453,0.00181868228948145,-0.0108699064332264,-0.0296447672032988,-0.00241369735384378,0.00747162273480795
"156",0.00751544756058165,-0.00290345849685891,0.00219454294321286,-0.0170048850285119,0.0103182337026178,0.00387091712860799,0.0257875096607931,-0.0218712845154195,-0.0219264640220684,-0.0171741360556121
"157",0.0183675041338811,0.0186921664566109,-0.00729928810442637,0.0316451724158264,-0.0040165207919769,0.000723002420348617,0.0262824826353094,0.0216508346031246,0.00510207173778587,-0.000794281750049253
"158",-0.00048389114647851,-0.00138272763484171,-0.0110294840483774,0.00204524165095177,0.000576397738478951,0.00216823166639224,0.0167010880156249,0.000520898865352892,0.00169206270751987,0.00278215339106791
"159",0.00200504599721785,-0.00277043551796652,0.0126393287714133,-0.00367351937541505,0.00483492484279391,0.00432615983454054,0.0150583958388728,0.011111167321687,-0.000767859301235019,-0.0015852880109033
"160",0.011867890372862,0.0247224519941809,0.0132162028047402,0.0430152974192184,-0.00160347372608327,-0.00323067636015928,0.00809158314394098,0.0317651409916049,0.00507149223912728,0.00238181403621773
"161",-0.000886204515056499,-0.000813364266582739,0.00724630508698665,0.00510574975833911,0.00344277031330931,0.000359937574004876,-0.00709021937604692,0.00931914671507617,-0.00137620790898463,0.00316823425738266
"162",0.0123534510600272,0.0215227529857969,0.00503587786601112,0.0238376439223793,0.00492033648111878,0.000359676628826522,-0.00633247933375092,0.0189611696989676,0.0122493190093194,0.0118436731577627
"163",-0.00930402573670652,-0.00894099627215661,-0.0078739609280396,0.00457994684368623,0.00523586994112168,0.00275904766015378,-0.0135590780128417,-0.00728132388911928,-0.0019663893213373,0.00117050424605614
"164",-0.0219803378497547,-0.0241178535339428,-0.00937946155824454,-0.0406535234598203,0.00169808757920253,0.0051438958951362,-0.0316155853395069,-0.0221676075186861,-0.00591098790947309,-0.0105221384053501
"165",0.0196216143952954,0.0259037942439122,0.00946826882168073,0.0396041688878754,-0.00271276987345648,-0.00380731661008393,0.0262600572817862,0.0218365809877881,0.00731825017949372,0.00945246275909684
"166",-0.00266161173504142,-0.0056212086793016,-0.00649368490666191,-0.00510437949228726,0.00668812056979129,0.00501739741957286,0.00484048038353135,-0.00897206560147068,-0.00408652943847421,0.00195096581230558
"167",0.00985283617629018,0.0171378171298595,0.0217863715832862,0.0258074331767095,0.000787968196491518,0.000237586743655704,0.0199589345194675,0.0139920764124721,0.0109421575558286,0.000389366640277888
"168",0.0100960034959887,0.00961550797941313,-0.00568552075851847,0.0168718028827097,0.000474065863094841,-0.00186093070617022,0.0134952180020009,0.0159086829516757,0.0138305027283752,0.0112884887874316
"169",-0.00865348757493034,-0.0139800689300233,-0.0192995932666494,-0.0151236413858125,0.00801740696214504,0.00621583027854555,-0.0239678860039801,-0.0209332132493349,0.0017793000658568,0.00192459985923144
"170",0.00230107941722735,0.00221555140549534,0.000728966992237678,0.00782713858132955,-0.00257672782050211,-0.00213816751411722,0.00613922795542821,-0.00522268211888599,0.01924220009598,-0.00384172346283407
"171",-0.0139068390101847,-0.0115826532923822,-0.00509856336470405,-0.0225592801875587,0.0141509365945576,0.0107142486619243,-0.0187122128056756,-0.0164071291810588,0.00769674691117128,0.00655603403984628
"172",-0.00191730260901746,-0.00581455922404506,-0.00878455482549201,0.000756844524342215,0.00775281682785378,0.00223909838881586,-0.0189304413844662,-0.0145121447972955,0.00331465633830019,0.00689651548866221
"173",0.0116609138825596,0.0197050166967021,0.0103398803051493,0.0201886583147695,-0.000769521643154913,-0.00211553854986868,0.018028348145013,0.0189572949562034,0.0129272329965284,0.00228314746503155
"174",0.00257681609210891,0.0032648055133746,-0.00292419264096055,0.00355800918959215,-0.00373900853440656,-0.00247320553463759,0.00179864551874376,0.010133175769822,-0.000850794137158162,0.0106301868737808
"175",0.00703279305797233,0.00562862121543861,-0.00733130684847505,0.011078410404276,-0.00894203225141532,-0.0059036283381696,0.0183678804679785,0.00970224314470558,-0.00539308835357777,-0.0075131534517725
"176",-0.0000674170681435049,-0.0099702948920718,0.00295424829890067,0.00197197858720921,0.00144801841231379,0.00130555932050536,0.00474579453490831,-0.00716630859494305,-0.00128430361631549,0.000757043374380428
"177",-0.00537230889982854,-0.0167841200482918,-0.00515463327301546,-0.00634234964657454,0.00478368783179994,0.000593629922908123,-0.00188924222004438,-0.0247704165006143,0.0140020435491368,0.0117245866427997
"178",0.0294396599715692,0.0420485978836016,0.0103626823733904,0.0484226914795836,-0.0075285329216922,-0.00106758629403947,0.0311022210890661,0.0277551882568448,0.0102859798466115,0.00373824050057459
"179",0.00590286007026841,0.00353470064488226,0.0109890590984605,0.00454836983919282,-0.00925643659468334,-0.00355994266480664,0.0203277445285879,0.019311927938811,-0.00376564869312324,0.0085661949880711
"180",-0.00704198024564262,0.0022338766914447,-0.00362306416853042,-0.0031347311915243,-0.0189128423374862,-0.0113150402537091,-0.012210815907076,-0.00851010557649778,0.0180596528069437,0.0155096524025742
"181",0.00269842064184855,0.00642977559066926,0.00218150805111983,0.0132776673016606,0.00849070209775515,0.00506001937126199,0.000260023399037523,0.0131573191312218,-0.00522559123727184,0.00690905679580123
"182",-0.00184222089381425,-0.00170349933992853,0.00362850028397355,0.0124139087060813,0.00284529374917253,0.00131838437577292,0.0085860133040665,-0.00145225099376101,-0.000829375218654893,-0.00180574604944927
"183",-0.0019782718207827,-0.00392524837151398,0.00578460217340471,-0.00374675109116029,-0.00351712066394461,0.000119437116717247,-0.0165533067508893,0.00226216399685186,0.000691795803704931,-0.0072358181019565
"184",0.00528462599401025,0.00436890398461842,0.00862667071467205,0.0133335159140298,0.000910679036156603,0.000358807162041508,0.00569005879926232,0.0169243671529911,-0.00456244975632647,0.00145768792851686
"185",0.00591355901618074,0.0119402320091639,0.0228085047827999,0.0148446097940229,0.00693866101452212,0.00323024351239676,0.00947355253332693,0.0112533513357602,0.0097221805555554,0.0262008927706412
"186",-0.00333128048862186,0.00463553919553861,-0.00069687848834965,-0.00631665379914459,0.00225952720178535,0.000358580665874797,-0.00325852490283485,0.00705379003384055,0.011141747364859,-0.00319145367419116
"187",0.0112729495561463,0.0100670261063789,0.0111575125399204,0.03144861105368,0.0057139965686146,0.0011959025681294,0.0265463255016178,0.00498030117976755,0.00530540048142014,-0.0103167347210077
"188",-0.00136092543701316,-0.00299013800754522,-0.00275865685635202,0.00681179384911523,0.00315048387977623,0.00215155372725362,0.00917210300103344,-0.00263242706736144,-0.020974343140072,-0.0201293040553866
"189",-0.00201205090662882,-0.0036653071966819,0.000691640551272243,-0.0302837427053154,-0.00291611211629017,-0.000715434191185693,-0.000252492515415592,0.00155264126077359,-0.00621970991623244,0.00110047505025279
"190",0.00156109705313012,0.00526756923347849,-0.000691162515249144,0.00996699379926258,0.00382509362817141,0.00178989033089039,0.000378707958136548,-0.00465118684690902,0.0134909731991384,0.013924485602435
"191",0.0118812817563922,0.00756869085074019,0.0131397788432843,0.0333551752787224,-0.0107577541520962,-0.00881527579955976,0.0198158242275315,0.00934563024348778,0.0072732122708985,0.0028913363212475
"192",-0.00532553405861136,-0.011474390079083,-0.00546082219599131,-0.0106321697025316,-0.000793061119841454,0.00360581839551322,-0.0111382882781348,-0.00925909813592118,-0.0118529015843896,-0.0209009532259744
"193",0.00941786894153251,0.0125262560312283,-0.00274531955252999,0.0155725477185169,-0.00124716375111555,-0.003113886349982,0.0057568364195355,0.017133751673323,0.00772090180230101,0.00699301195640767
"194",-0.00166154393399387,0.00041245630274056,-0.00206471551512133,0.00133068296675587,0.000567570166956743,0.000961696733222883,-0.00136904999318621,-0.0013781899491172,0.00369414440794325,0.0116958755188288
"195",-0.00480049574069563,0.00412195715604646,0.00137948613179595,-0.0087954902821622,-0.00102096340275959,0.00011924461495938,-0.006728822645649,-0.00398713182626254,0.00749731451066915,0.0111994302013048
"196",0.00553096896719407,0.00615771295669698,0,0.0182581608344197,-0.00488295307390729,-0.00335974401577699,-0.00727628722141205,0.000770197507512282,0.00920027010146018,0.00464463410506832
"197",-0.00844347932800471,-0.00873119834018177,-0.0117080616789698,-0.0122254824857729,0.000228396669471609,0.000962947840107198,-0.020598950329254,-0.00846175061042109,0.00737368319472775,0.0170696735864164
"198",-0.00793493710556148,-0.0113599583306038,-0.0181186282276603,-0.0185340207238018,0.000342474845667073,0.00276646543273062,-0.0166454605730256,-0.02172244860672,-0.000266116585921239,0.00104887679717081
"199",0.00305626094177058,0.0122396197606995,0.0014196274065017,0.0230872795735688,0.0109484517598613,0.00611821634719423,-0.00275533549165696,0.00475852533797938,-0.00825350073535003,-0.00523930066369616
"200",-0.00363018308698049,-0.000493161428931188,0.00425211008107773,0.00505718235900465,0.00552785436926384,0.00381559183401858,0.00263163877436634,-0.00552551555269976,0.0201342281879195,0.0179073168434274
"201",-0.0261567457504568,-0.0198337524712986,-0.019759994230043,-0.0427675581404313,0.0149224216159303,0.00855216656844404,-0.0322832457820391,-0.0273012911263851,-0.00394740789473691,-0.00275953735000611
"202",0.00581265277407228,-0.00503802543375953,0.00575952700521576,0.00722743274676785,0.000109853769357349,-0.00188439627053039,0.012340358367334,-0.000489405935752529,-0.0145310309589576,-0.00276717346854638
"203",0.00810484024939062,0.0156116832526456,0.00286331605762569,0.0277236218169916,-0.00132640355679137,-0.000236292812642702,0.00870729750144461,0.0179593828917843,0.00844510746501625,-0.00693725997684724
"204",-0.00184568155914056,-0.00124617849323672,-0.00428287454962073,-0.00653767605790867,0.007415831955492,0.00507519463087669,-0.00398422087581429,-0.000160481676568902,0.00385476523243011,0.00349284216203993
"205",0.00237703363350006,0.00582366948441537,-0.00358395473917084,0.0127139193431693,-0.00340609348923626,-0.000822133854137763,-0.00266681677694236,0.0131536296805252,0.0067532047174208,0.0233204754837524
"206",0.011722580365066,0.0168733686694333,0.0172661709227624,0.0283262004676803,-0.00231416947206309,-0.00246780824299675,0.0147062213875242,0.0186826168858916,0.0218335265268121,0.0153063169226604
"207",0.0033199804375128,0.00618192787911753,0.0134369908488996,0.0230064055465338,0.00386670221149599,0.000825326060855947,-0.00724645347326114,0.00326400027556017,0.00553483059506155,0.0164152409450689
"208",-0.00694244809718925,-0.00727582582120334,-0.0048848306186946,-0.0188906239391676,-0.000550276837403274,0.00105910238470042,0.00451223269080647,-0.00325338123830199,-0.00985669444994774,-0.0224126033472398
"209",0.0103878825808537,0.0146580370246554,0.00701270386690056,0.0219437450420219,-0.00903018559305802,-0.00670283111559145,0.0179679879503227,0.0219146810515911,0.016418940308182,0.0283210275855652
"210",-0.0234070848166953,-0.0244780525440389,-0.0125349077734968,-0.0403734296779785,0.0129926334228718,0.00816175276716713,-0.035691146280739,-0.0267679887188113,-0.00877643059871147,-0.0127869289061899
"211",0.00112531797239557,0.00822698204061978,-0.00282082543272433,0.00567216104827173,0.00319563953400226,0.00270977469542699,-0.0197845080661635,-0.00781355895308733,0.0243808802771717,0.0215875633978628
"212",-0.00760577024457576,-0.0134639589602653,-0.0169731102992449,-0.0347693525705844,-0.000439269567567013,-0.00117467460733767,-0.0142796138821086,-0.019530589363744,-0.00100215455337194,-0.00650202454672566
"213",0.0134621309907494,0.014061189658737,0.0115107879267731,0.0379477957054286,-0.00483543971624523,-0.00176510360746718,0.0104470242287529,0.00883506238237364,0.0210658307210032,0.0261779946862162
"214",-0.0273561102043502,-0.0160685751616176,-0.0184921031570132,-0.0318586007506626,0.00176692505198761,0.00365437467862773,-0.0337749583881595,-0.0195854770303301,0.00994716934790607,-0.00510201048791581
"215",-0.00507059572953239,0.00887016921766315,-0.0159420700350371,0.00511174065717657,-0.0017638085345012,0.00223110226869294,0.00627810760800918,-0.00357370777433452,-0.000121534536029588,-0.00256400139839019
"216",-0.0137259744223902,-0.0230074636117131,-0.0132550599377554,-0.0235220793747982,0.00850308741987305,0.0059757145043644,-0.00340303605273573,-0.0203748910244881,-0.000608087050659512,-0.0003214058130524
"217",-0.00992183156022874,-0.0159797958228595,0.000746193248328808,-0.055338617748541,0.00361366770798388,0.00174791126653706,0.000142617758093433,-0.025790174044641,-0.047213397420297,-0.0218579729895122
"218",0.0304800078146155,0.0286323042383279,0.0171516258180291,0.070640893701329,-0.0037101138569503,-0.00511621888344926,0.035846308333239,0.0401367657881879,0.0104725411057773,-0.0190600112852922
"219",-0.00276865385461234,-0.002907922456026,0.0029327686213807,0.00096552479408718,0.00109522358084835,0.000701090714426256,-0.0146938047534559,-0.010673523748897,0.0146612229021277,0.0224454312693505
"220",-0.0144239819123486,-0.0166668674288888,-0.00877206530936858,-0.0230222564211353,0.00940774413587131,0.00560549197423121,-0.00557478342616102,-0.0182571756651423,-0.0290234433112039,-0.00982962716745794
"221",0.0017175200138817,0.00423735890730281,-0.00737489607814812,0.0123747487973558,0.00140861607570453,0,-0.0190609430765264,-0.00422645500607266,-0.00256570888642882,0.00330906930670882
"222",-0.0139242384306673,-0.0270040373328425,-0.017087458515992,-0.0460988745753405,0.00649194192699265,0.0072017156024331,-0.0191456992002431,-0.0280136611548559,-0.00655951125401932,0.00758579294261863
"223",0.00612146709106187,0.0222893732384184,0.0264551136382229,0.0274694643217368,-0.00107478848530196,-0.00265332423622167,-0.0233064502695743,0.0155455561737017,0.0288710908563203,0.0248772327886559
"224",-0.0204643522986581,-0.0184947107678094,-0.0176733683470071,-0.0503518073806842,0.00581196442787713,0.00786315700630569,-0.00745726412202941,-0.0223592629369876,-0.00138417010967451,0.00127765068033292
"225",0.0172923226803314,0.0215228047988809,0.0224889755431115,0.0295495104461703,0.00299674729300659,-0.00298301490848951,0.0190835312523492,0.036241876792906,0.0238155112926473,0.00925023354463761
"226",-0.0220635262222151,-0.0197156590077066,0,-0.0396933255160701,0.0197373920182087,0.0136925763127711,-0.0376001268154023,-0.0290319248164166,0.000615421538461502,-0.0123260774232595
"227",0.0114935938318159,0.0125163116857656,0.0161290762428195,0.038295627060162,-0.0095212568228058,-0.00930736428996948,0.00735438587086268,0.0307738637235435,-0.014760208557434,-0.00800003976861519
"228",0.0319841116838209,0.032395627971058,0.00937954955064146,0.0547809002287301,-0.00676039944433393,-0.00355225777096235,0.0468442034314593,0.0154373621997981,-0.00661670428506134,-0.0122580734124823
"229",0.000339684599770518,-0.00908339034742622,0.00357412063628049,-0.0122583817324197,0.00861466138759703,0.0056337839177405,0.00799076170573443,0.00133618249152168,-0.016212152821415,0.00228622915887211
"230",0.0100561297776358,0.00374993324759165,0.00213627480086309,0.00849140201305798,-0.00484998147134441,0.00137218570626341,0.00922420122686352,0.00600611586476307,-0.0122636562629492,-0.0123820652419223
"231",-0.00659253283735517,-0.00356973706323627,0.00142166731415938,-0.00867886485765412,0.00793494931996319,0.00395276358858987,-0.00728309967593077,0.00364855558623334,0.0124159208484222,0.00725844226775885
"232",-0.00893843819084317,-0.00599911014930588,-0.0106458314714766,-0.00261346672342477,-0.000105404799972342,0.000912752726109689,-0.0261835631471921,-0.0133845370084552,0.0143076522011707,0.00458558632946859
"233",0.0167398707445374,0.00813033636826654,0.0186514443211649,0.0444125040982775,-0.0119271387255083,-0.00376190226834938,0.0285120416011642,0.021772236913413,-0.00969779572549634,-0.00749915544072055
"234",0.0143134926349608,0.0106432339443117,0.0126760610556844,0.0157425812077283,-0.00875956757919738,-0.0052648401091081,0.0359097841572571,0.0136043517195499,0.00941124288736761,0.0180682734706157
"235",-0.000198134643352832,-0.00255058005367281,-0.0090404572675431,-0.0118554288381991,-0.0112084126218612,-0.00644198818835862,-0.00485322438230229,0.00258721156381436,-0.00970146114269388,-0.00322681525340973
"236",0.00775253585854396,0.0112174403718421,0.0028070545852994,0.0003123725231029,-0.00599414335463511,-0.00231628127598416,0.0250800344230475,0.00403252082865468,0.0178117307331229,-0.000647459196076228
"237",-0.0274200709629402,-0.0268354472793245,-0.0216934520423043,-0.0423538026959146,0.0196267098043605,0.0136953350995945,-0.057224321012054,-0.0224901784847698,-0.01450005,0.00874629264896143
"238",0.00987127052225056,0.0233846377821265,0.00786832850726782,0.0300065800351814,-0.0103236541926136,-0.00835783609912877,0.00317178924963146,0,0.0209284891389392,0.0272961382131933
"239",-0.00207589047483026,-0.0197377474614493,-0.0205817735031592,-0.0274857963272479,-0.0108659151225062,-0.00739008649775386,-0.0172466551069168,-0.0164340263431867,-0.0247235439116299,-0.0106282956909713
"240",-0.0126793511457917,-0.0252319824711406,-0.0391302905008757,-0.0238343651268929,-0.00461318098470909,-0.00290753919575715,-0.0302717110990147,-0.0342517244055561,0.000254738853503245,-0.00695106564738879
"241",-0.0142690497171404,-0.0173996515001944,-0.0173456162983323,-0.0426284500170245,0.0089382670469953,0.00594930117621795,-0.0180969526305428,-0.0501731653601776,-0.0049668876069876,-0.00489079563714301
"242",0.00558365400895222,0.0109911334849944,0.017651797606592,0.0274541672722677,0.0064541627801602,0.00197148163678973,0.0129010110658769,0.00273182780341674,0.0143351215026926,-0.00425944207669848
"243",0,-0.0101812337251252,-0.00678758402537016,0.00651120818455642,0.0132595635737063,0.00798662826711882,0.00834004648687436,0.00999085374572761,-0.000126208201892797,0.00954259968372395
"244",0.00630688270873514,0.00392273149096334,0.00379656263773898,0.00545770162214598,-0.00214496672721609,-0.0016075306303065,0.00375950900778732,-0.00629497538809787,-0.00719333688019519,-0.00423733058600284
"245",0.0144150289937499,0.0145870394909495,0.0151284440555808,0.0301568659019555,-0.0146191483949967,-0.00724564388029714,0.0170785976426768,0.0130327279147264,0.0181771963436428,0.0117839818799261
"246",0.00742578804651073,0.00679760470341573,-0.0016561270464257,0.0169132388094759,-0.00469003051782191,-0.00289670187424984,0.0272501872729904,0.0189188322507157,0.000499388277138246,0.00744093606279606
"247",0.00214413199888219,0.00550257946184884,0.00452475929424789,0.00518333649456926,-0.00876860601275198,-0.00476372553720994,-0.0166332855484492,0.0150307041861906,0.0172198404943829,0.011881835103565
"248",-0.0125706913420595,-0.00277981780909575,-0.0157657196913448,-0.0230757794527133,0.0109021223220855,0.00671393459252334,-0.0194549395030403,-0.0243897581012811,0.000490689419431423,0.0034910490379898
"249",-0.00250576557609516,0.0083624485930256,0.0114417287112698,0.00376082974259884,0.0155933503178141,0.00803155085487672,-0.0147412473634319,0.0157141080076471,0.0176557385398661,-0.00316255885803629
"250",-0.00739962455731569,-0.0122668470739286,0.00226229999748773,-0.0120290131569113,0.00605568791236877,0.00461760087716279,0.00305362818437849,0.00123075516631155,-0.00650603614457834,0.00126896397825904
"251",-0.00875487358518101,-0.00271119474158721,-0.00451475038780724,-0.0165006262338848,0.0144020156882563,0.00712591106770666,-0.00837176835988274,-0.0043897481982742,0.0291050452231998,0.0275666024282257
"252",-0.000482679995943647,0.00175388613183647,0.0037795525084825,0.00899752046815827,-0.00137768108339764,0.00205375240091277,-0.0323865701478838,-0.00370391814164173,0.00836670977649412,0.00770883958221713
"253",-0.0245065507350612,-0.0234611337288972,-0.0256027168065389,-0.0300367093628903,0.000212496929970829,0.00261965763766714,-0.0317256677248479,-0.0219507017469422,-0.00514202407385755,-0.00581387407030654
"254",-0.000849284816573537,0.00502004387097243,-0.00618240969955097,0.00732701731362817,0.0043493781149373,0.00181770926549496,0.00933815771063329,-0.0162893925341892,-0.00422882664967084,-0.0181595601336975
"255",-0.0161483497168555,-0.0090983756862919,-0.00233257387666974,-0.00775398419664874,-0.00116271922918409,0.00215386358120173,-0.036358050972654,-0.0220791375625529,0.0237112430238733,0.00909093024415042
"256",0.0105101154725269,0.00414108391558377,0.0218238322022217,0.032780035162097,0.00190400604462337,-0.0015836672297902,0.0197072508136877,0.00564456273892677,-0.00265033420892291,-0.00994093566611409
"257",0.00655406359196542,0.00080654537714353,-0.00839049364031019,0.0117850873317003,-0.0135094003344834,-0.00271979327602967,0.0132142813915139,0.00187035695232951,0.0196417901915036,-0.00470664262171938
"258",-0.00806853492951176,-0.0173774248952824,-0.016923188341543,-0.0281268698933901,0.00781064094608341,0.00636328802849628,-0.00162994336807087,-0.0252097613376174,0.0037393994334276,0.00914241888765055
"259",0.00806303810587128,0.0165908766911871,0.0125194310083654,0.0147085456828111,0.00371513424135328,0.000451506759426623,-0.00277629797185264,0.0153255008208799,0.0108376493376012,0.0124962089895626
"260",-0.0220131592534148,-0.0312948853451521,-0.0278207503687156,-0.0452318519054824,0.0112107363021445,0.00654465955419292,-0.0260355192370284,-0.0309433854830699,-0.0173107324401304,-0.0123419810154484
"261",-0.00861244151085194,-0.0216602871597643,-0.0182827229913249,-0.0416109231734758,-0.00721652056745259,-0.00190572093248786,0.0129455362353013,0.00272606517712393,-0.0146607686023587,-0.00937191995711351
"262",-0.0259162609892999,-0.0142874774960327,-0.0137652874200634,-0.0291160514565815,0.0129579250188132,0.00808858111873678,-0.0121161379726323,-0.0108742401678492,-0.002306770552714,-0.0129297788189532
"263",-0.0102677125646341,0.00105619261927825,0.0262725761660576,0.0228130963657633,-0.00686377111050263,-0.00144885374167747,-0.00840063585598916,0.0070674630866856,0.0106358150289019,0.00383388391305206
"264",-0.010146520057257,-0.0312591271691831,-0.0368001830828457,-0.0251110742622984,0.0106813725931441,0.0111596406660306,0.0337170919486358,-0.0183234353779052,0.00857927267397107,-0.00350091581404965
"265",0.024020966878314,-0.00653265262722247,0.00332235039548401,0.00636346992283299,-0.00227938901686886,-0.0046352811027135,0.0817901909583658,0.0127082112432764,-0.00317567206931324,-0.0188438187034397
"266",0.00844154521581086,0.0297896072831794,0.0165562700501978,0.019421961299356,-0.0200435978070336,-0.00909196847251093,-0.0195456882447534,0.0284314787191773,0.0249175449416035,0.0247395512072714
"267",-0.014445658297552,-0.0201239640770395,0.0154723926063782,-0.015211690906119,0.0168509723900396,0.0092871706444293,-0.0139078985872768,0.0285988913321134,0.00244228458165452,0.0222363674138357
"268",0.0165364786057491,0.0156991348390574,-0.00561323851586082,0.0247448081112029,-0.00375301122568261,-0.00365911313189426,0.0371413128569904,-0.00185377598344083,0.0160575520689628,0.00466139951663203
"269",0.00495400481560826,0.00767967676365577,0.0169351638415072,-0.00490249583913993,-0.00679980054918838,-0.00400559155612212,-0.00604420398035066,0.00185721885114321,-0.00653948773841961,0.0083512203980638
"270",-0.00735762638942583,-0.00347268800631062,-0.00475801954107113,-0.0131627287772461,-0.00652981849102163,-0.000446990819266246,-0.0234114168846141,-0.0157556795039731,0.00998349950667032,-0.00858889055647272
"271",0.0182341912196182,0.00948668547636156,0.0135459459602427,0.0200448985139179,0.0071031078292263,0.00514164136900819,0.023817119665718,0.0169488734431582,-0.00716919415966089,0.0049505395663092
"272",0.0160878798822113,0.0138090510612461,0.00864777268771433,0.0199425906083033,0.00601141231062008,0.00324630430043871,0.0389235549595028,0.020370840592453,-0.0224289272991482,-0.0175493094837592
"273",-0.0126091355113472,-0.00813448715664822,-0.00311789527239914,0.00308002919000505,-0.0102917111695822,-0.00555919313949571,-0.0155134723270287,-0.0038111572010624,-0.00279798551310539,0.0175493516543039
"274",-0.0267738186921639,-0.0500670187854794,-0.0336201815651371,-0.0538380055091345,0.00763999025414397,0.00704380200488397,-0.0316631394517809,-0.04354150680277,-0.0159371271815292,-0.00831537447744168
"275",-0.00805193572777951,0.0055215656334151,-0.0129448523459926,-0.0163761735563973,-0.00305398714319483,-0.00177618905030341,-0.0191893269192912,0,0.0144844548357663,-0.00465840677163776
"276",0.00661376202714936,-0.0108826771651727,0.00573776336801601,0.0169557751738949,-0.0215457257763844,-0.0112333315566221,0.0241040515374531,-0.00857159712211242,0.0101180554283773,0.0121684457745848
"277",-0.00642109009592884,-0.00353272758099421,-0.0252649012151912,-0.00188632406186073,0.0114413165359948,0.00843612713892283,-0.0310254853263879,0.00192122226798186,0.0127991321713774,0.0299014221653737
"278",0.00510970275880451,0.000911718154646524,0.0100334674308051,0.0123962256642085,0.00416299660523212,0.00223043975949322,-0.0200315682905591,0,0.00362639560439559,0.00658490632753428
"279",0.00927147222701619,0.0254022453868097,0.0149005955831762,0.0161266869160333,-0.00595239468252873,-0.00211452135748003,0.0315466066780221,0.0134227677555627,-0.0218986089587516,-0.0202200517606466
"280",0.0102228983130694,0.0141137162590976,-0.00734087688391361,0.0224835215121146,-0.010584005946857,-0.00423813858684952,0.00468071061823983,0.00851461389634856,0.00123138920337218,0.00819414455935585
"281",-0.00879980255674517,-0.00778599842136729,0.00986025982068672,-0.0128629709769462,-0.0146968842190807,-0.00548772677778375,-0.00745445086771268,-0.000938137272696871,0.00301874993249651,0.0201685945015921
"282",-0.000221749127788384,-0.00392306628506423,0.0122050357416772,0.0071343357271676,0.00767779199652829,0.00213943126359184,-0.00406817061851639,-0.00187770944514343,-0.00624230304583995,-0.00472116848927839
"283",0.00281178534400373,0.0125059915315988,0.00964661540929423,0.0130824798197509,-0.0101226955606952,-0.00719215089654657,-0.0174393613563928,0.016932960280599,0.0272574306840732,0.0326120194826895
"284",0.00295166260544932,-0.00048654988345731,-0.0207010302620606,0.00834791206910324,0.00692684712171454,-0.00090634318717786,0.0233454062776672,-0.0129512463919329,0.0181261843606424,0.00516786232688937
"285",-0.00831389162205698,-0.00136201347290987,0.00731734818200858,-0.0140099456669825,0.0105917970012088,0.0103110745967363,-0.0226564336513827,-0.00674744077845535,0.000107271559572464,-0.00542700647917216
"286",0.00615774797579216,0.00964653537819626,0.00807102578679952,0.0134194314657685,-0.00572610752680902,-0.00280383842206677,0.0235012980625828,0.00490642874027203,0.0015013297587132,0.0137852753837973
"287",0.0126086476119849,0.0147652699882279,0.0208167857480752,0.01862334506972,-0.0102152728891295,-0.00663540297176946,0.030928016035294,0.0140841468276003,-0.0069600707459051,0.0096317030604518
"288",0.00750073902819981,0.0194958227338011,0.01098038230012,0.0132081545501372,0.000329252614199138,0.00248983329702179,-0.000606283791675821,0.0138895416802678,0.0104593597252396,0.0213242670851113
"289",-0.00101212056875688,-0.00335833460404167,-0.00543087754719218,0.00843902086719939,0.00087755387926558,0.00237257925603362,-0.0071253664310994,0.010045675523829,0.0114182052226892,-0.00137369983327418
"290",-0.00976722396386298,-0.00393130458355961,-0.0109203599239003,-0.0107494696568509,0.0177650756501286,0.0117174119619337,-0.0207667689763165,-0.00542507327450281,0.0127663959988014,0.0096287237141659
"291",-0.0222836538594927,-0.0247131485550178,-0.0118296197772652,-0.0397527764928246,0.0153007169824375,0.0106896491721176,-0.0174643480822699,-0.0334546563695965,0.00197939372808409,-0.0163487644500253
"292",-0.00239147143978369,0,-0.00079805824611423,0.00544369740651884,-0.0025779837275306,-0.00254145915922865,0.00539591367051484,0.00169293409802229,0.0110209814930338,0.0146813734667879
"293",-0.0038201125315156,-0.0112725307564474,-0.0231630174749682,-0.0232226880063058,-0.00971793860842807,-0.00376758112125786,-0.00805018358513876,-0.0159622558858745,-0.0211846775233376,-0.0035489822077398
"294",0.00631611576003555,0.0109138890969507,0.00572349109072445,0.0210033438310371,-0.0119700024964807,-0.00433688433324741,-0.000955052269841383,0.0160306869257536,0.0266862891363731,0.0219177486587276
"295",-0.0206979401160468,-0.011374833244097,-0.00894296760257418,-0.0342856839223376,0.0053475357793098,0.00804202740743065,-0.0458746346124095,-0.0159655029966975,-0.0124846601260268,0.00750686883795959
"296",-0.0103002933302854,-0.00887259595378231,-0.0147660370923232,-0.0138316879358137,0.00130298349195868,0.00343570219924816,0.0100169968268367,-0.0112619165101455,-0.00424874611398962,-0.0101118449885799
"297",-0.0131832823562256,-0.0102313469504068,-0.00416336097617542,-0.0175500537545958,0.0147454916592205,0.0071781223096945,-0.0161983101526281,-0.0173738556114779,-0.00228944748837334,0.0188172265118327
"298",0.0359375906360933,0.031806265514988,0.0292644355954432,0.0672569594401005,-0.0085474041497986,-0.0108554173400141,0.0710679424823726,0.0451863289592842,0.00125164281052537,0.0155672258795234
"299",-0.00935165284306805,0.00250418363338079,0,-0.0185264349540042,0.0192904633825357,0.0115285446014952,-0.0214895125194619,-0.0203007637453879,0.0106261487785426,0.0109120036113952
"300",0.00220778241340835,0.00490082020347637,0.0032494055348169,-0.00910989375559546,-0.00782406659510115,-0.00525964287259451,0.0125035564308817,-0.00230275578351102,0.0137098646797265,0.00102792855388745
"301",-0.0154960052246771,-0.0253393864126886,-0.0663968792273657,-0.0354518500479746,0.0123620251062517,0.0103550259497138,-0.0163075669163257,-0.00576898631083633,0.00376248744203722,-0.00128365835410771
"302",-0.0101070564544704,-0.0171690388768914,0.0286210895299339,-0.0247063680755417,0.0076836618905316,0.00501664109214217,-0.00676001181100816,-0.034816372717685,0.00466010540634287,-0.0401027999348437
"303",0.0415434021621297,0.0303457191261616,0.0286675528931388,0.051993507098774,-0.00386422504536865,-0.00683619951336945,0.0510449538503777,0.0320642002752094,-0.0269234451330734,0.0222280619906789
"304",-0.0247699129477563,-0.0382679230349828,-0.0303275877127035,-0.0600519033094605,0.0165685001116158,0.00863120742388457,-0.0109464006314234,-0.0194174757281553,-0.0358549119170984,-0.0432275970356528
"305",0.0185227492741316,0.0126927838375328,0.0185964252834616,0.0168424093909199,0.00247578212819866,0.00216520886894656,0.0417767499011903,0.00406200850057226,-0.0336414119342067,-0.0402519045767038
"306",0.0199878607655057,0.0179050834557806,0.0307055873794548,0.0383354698969915,-0.0193461486754267,-0.0176159732472809,0.0170581477588825,0.0392706831703584,0.00211315750803442,0.0182596148216252
"307",0.000965147423514168,0.0177855809852951,0.0104670073118829,0.0153525524083113,0.00419777366065843,0.0035209741447535,0.00788450428135756,0.0095421757796581,0.0291898452650354,0.0100869355330777
"308",-0.0122358143630206,0.00384050258767243,-0.00796820067726134,-0.00811343802672027,-0.00418022601798451,0.000767651218092302,-0.0264204945964733,-0.00378085877111589,0.0115388759342541,0.0299583839720059
"309",-0.00315357614037992,0.00124378250344637,-0.00321303627346925,-0.00483329928329834,-0.00702970378053613,-0.00131516060586312,-0.00424503560785472,0,-0.00362477600347211,0.011042175200366
"310",-0.00956448580254288,-0.00487234229195932,0.00402916849348856,-0.00179380326122958,0.00972180499233777,0.00394924150530618,-0.0153775602522174,-0.0153700536687479,-0.0169056496565979,-0.0237079151963853
"311",0.00349788587233602,0.00806374909955876,-0.00722292432046645,0.00591409148514632,0.00355864654085725,0.00174693052674635,0.00664912847719856,0.0185005494098731,-0.0159990536351454,-0.0240109860613007
"312",0.035159453704251,0.0318065186247996,0.0291025079486005,0.0383985241808344,-0.0162749517763143,-0.00874317091172838,0.0491551897948201,0.0454115682018492,-0.0392655994130915,-0.00559131338682139
"313",0.000658780392421177,0.000369075267574459,-0.00157096895453568,0.000716633334819416,0.00212922312743324,-0.00331181393409885,0.00424601392392221,-0.00271512946217323,0.0277457514650501,0.0298003766841444
"314",0.00248741648349093,0.0016609188491743,0.00472058350334259,0.0121742355850873,0.00223069928310471,0,0.0204114898210015,-0.00181430444418884,0.00168030699048871,0.0054601548488511
"315",-0.00109478989389489,0.00543389247927939,0.000783154026538169,-0.00403298502223071,0.00911591121833744,0.00764257249270606,-0.016288302784385,0.00090871362706002,0.00928206238608942,0.00705930535222699
"316",0.00051136582575384,0.00494694799370965,0.00704225668044756,0.0132840658539539,-0.00525239497664032,-0.00659524707569159,-0.00232379821269091,0.00999051367864068,0.0101938836565099,0.0107847322711923
"317",-0.00102214346133411,-0.00911565161078509,-0.0147631125211509,-0.00546814508717575,-0.00348449996930522,0.000110280495087434,-0.0125199656062055,-0.0151078276237402,-0.0089941868815222,0.00400083423797892
"318",-0.00723582671554013,-0.00386374259821576,-0.0149841136572572,-0.0155787374285492,0.0103843371256149,0.00597493795951398,-0.0203450598299894,-0.0189915573601849,0.0214720868062444,0.0167376768781422
"319",0.00139894724660139,-0.00295541773186092,-0.00320267348738845,0.014321348574176,-0.00335565104733815,-0.00396008250425717,-0.0021066940701463,-0.00874924350914641,-0.00563445654313077,-0.0044422060963667
"320",-0.0194088843838197,-0.0163023374989669,0.00642573322021489,-0.0163073590625794,0.00673483523140761,0.00430718033940436,-0.00361992972805381,-0.0101408098010332,-0.00512143418725408,-0.00393697157603001
"321",-0.00337366830639085,0.00197738932821223,-0.00638470679764391,-0.00236877598460072,-0.00585401945594222,-0.00252879667080785,-0.00544826315259006,-0.0098652322484265,-0.00208107331606555,0.00685105097014449
"322",0.00233188987881627,0.00488694552752467,0.00722901652620522,0.0117260715031884,-0.01240590126509,-0.0045194964145282,0.00517413284795798,0.0136043800690142,0.00603669184461975,0.0120387266780331
"323",0.0270940183002377,0.030113234305936,0.0318977856301266,0.0295786229157433,-0.00979416964706903,-0.00675481611691253,0.0431492268879496,0.0302454520059843,0.0175648366762018,0.00956836643833903
"324",0.00146114434320221,-0.0128008677391658,-0.0146828790691477,-0.00725117863229463,-0.00172110021577065,-0.0023405966184995,0.00580542100027315,-0.00422050910614646,-0.00761229787538231,-0.00461070342382686
"325",0.0104344933756271,0.0121388559075113,0.0274508255800376,0.0150956974907941,-0.000861608608368369,-0.00100584031319428,0.00101038087449346,0.0068177812066692,-0.0209593241348168,0.000514571753596815
"326",0.000505290799910352,0.00254420062722249,-0.00305326500725045,0.00507091566223616,0.00398858512101508,0.00011111961689414,-0.00994705301399434,0.00311150562836038,-0.00408301685887158,0.00128607698844219
"327",-0.00440251043201267,-0.00879093676211029,-0.0191426380429406,-0.00927299782225044,0.00343516346836581,0.000783841616459169,-0.00465912449011541,-0.00437889214579712,0.000221573407202191,0.00616493979980648
"328",-0.00159511993737038,0.00128011234584346,0.0109291190492231,0.0143842765185924,-0.00331582939807484,-0.00100663715382121,0.0115563210473899,0.00293198328244992,-0.0116317274276636,-0.00944611904816373
"329",0.00435680313709108,-0.0039267186951355,-0.00772198451017303,-0.0128230846853411,-0.00848169258092901,-0.00783039793952334,0.0229934249572354,-0.00876998963189779,-0.0224164982916779,-0.0167525302708712
"330",0.00925389646555619,0.00980952519158862,0.0194551235325855,0.00735372538331847,-0.00584627769336477,-0.00135245735577549,0.00339298370829311,0.0046081921509149,0.000573217145457328,0.0183485356086419
"331",0.00021512255103695,0.000725956896574731,0.0183203271632113,-0.00191032624652776,0.00304972263061987,0.00180595414813012,0.00225381132452407,0.00642207342922063,0.00481270785422394,0.00231666710798772
"332",-0.00393900126536784,-0.00816463469936068,-0.00899518457732829,-0.0177045298650366,0.00379905470631292,0.0018032537738828,-0.0144780831692404,0.00182327480481748,-0.0214392058059254,-0.0241397522296555
"333",-0.00589617905128925,0.00301844962138209,0.0045387243295103,0.0205982040986064,0.00713944835566727,0.00314988650977899,-0.0175442872640281,0.00873459409025412,0.00978911571586338,-0.00184207728080377
"334",0.0206853723918363,0.00729540639032056,0.00903575308970539,0.0106372088748568,0.0000648117394719261,-0.000112541069389849,0.0235194403701804,0.0073969359631143,-0.0306982566486265,-0.0232005671045774
"335",0.00276384897593474,0.00153912990063376,-0.00223866480447166,0.00958044653984591,-0.012610985993987,-0.00810056871221176,0.00170190798996406,0.0109241097620298,0.00702469358315727,0.0253710588069842
"336",-0.00480558158898114,0.000632465966605045,0.00149592719826974,-0.000735286030412841,0,0.00147428994994336,-0.00240672229287375,0.00212595720551878,0.0199810234102384,0.0207949517827233
"337",0.0086633817696995,0.00505877370284136,0.00448067257820139,0.011168249595348,-0.00720417285406016,-0.00317121180817814,0.00794864386605454,0.00212103905070382,0.00417294554907666,0.013151143431118
"338",-0.0178108014685724,-0.0171670004509912,-0.0126389235985916,-0.0297617191848609,0.00428805070019411,0.0039768139958154,-0.0294324801321904,-0.0225788042891826,-0.00935007535553778,0.00178157001672608
"339",-0.0025803713101975,0.0075902576381297,0.00451760387166833,0.0102930032753616,0.0089774267788405,0.00645141035693797,-0.000435343580409753,0.00721901082211129,0.0165462363085529,0.016260283314486
"340",-0.00186815528028483,-0.00599032647688291,-0.015741725699203,-0.0081640275609236,0.00368993840087484,0.00112399341851388,-0.00711288739217542,-0.00662944490871697,0.00206327377494908,0.015499896788278
"341",0.0112312019605247,0.0114135023851376,0.00380815349198849,0.0128573156878955,-0.00151424261057753,-0.00168495444260108,0.0213453032887851,0.00270530339601649,-0.00491878299974347,-0.0169866569386756
"342",0.000142427497126452,-0.00496527201545183,0.000758516922436892,0.00476851142217694,-0.010935059173144,-0.00832569111832004,0.00529634483378483,-0.00845461705873529,-0.0183929076535903,0.00550965867879594
"343",0.0020639472037427,-0.00217740539100986,0.00909775205335239,0.00240609964695238,0.000437503591324662,-0.000340420779720407,0.00669206114149157,0.00598654211958372,-0.00222510835256018,-0.0161893475568939
"344",0.0125030203070735,0.0136387953676942,0.0195342197079971,0.0212723520185605,0.00908140902033905,0.00556119066190086,0.0124471460372209,0.0126244107789018,0.0211267965185493,0.0113924318653231
"345",0.000912198614168469,0.0123789875322151,0.00368443206703861,0.0127329966645875,-0.00412001667126538,-0.00169292239134233,-0.00656671554842314,0.00195910296338919,0.0241379080459769,0.0145181541236565
"346",0.00273380549787317,-0.00301269783930613,-0.0014682253796966,0.000193391853545721,0.00130722158515484,0.00226056244926998,0.00759441867895339,-0.0120872595947711,0.00325478121784029,0.00148039177348736
"347",-0.00810918589501175,-0.00684319591345428,-0.00882381420275491,-0.017340530896388,0.005218824898088,0.00304649242757016,-0.0206561166293897,-0.00791608953400302,0.0168923035786139,0.0137964968803499
"348",-0.0169146532722806,-0.00912729997061545,-0.0178039729590395,-0.0101679883212435,0.000217325217052977,-0.00236226587715405,-0.0216615214395164,-0.0126948925399362,0.0116611328567406,0.0291615105691487
"349",0.000143482225550384,0.010566024210211,0.0143504354072919,0.00291621808290232,-0.0117891798898774,-0.00653781572755241,-0.00670076904746397,0.0121231670837201,-0.0106567639262372,-0.0144037392189068
"350",-0.0134042753368706,-0.011974874380291,-0.00819050513908282,-0.0174453356779577,0.00437713032408737,0.00442479782002336,-0.00645288348600281,-0.00980039997856441,0.00274785658118737,0.00191664407877123
"351",0.00741055148548098,-0.00388913916796607,0.00300292626332488,-0.00161422063286132,-0.0067556430357999,-0.00485672157064443,0.0143175224519385,-0.00751439042097757,-0.0204976645676532,-0.0160210091301101
"352",0.00461567336157875,0.00381346745494704,-0.0112275129574287,0.0134727051604808,-0.00888600091169933,-0.00749288727853781,0.0040745660672048,0.00757128400497908,-0.00246197401004944,0.00631828367677323
"353",0.00502522479047407,-0.00597009473372501,0.0113550013825834,0.00219323937913174,-0.00719593248229144,-0.00468933903155155,0.0104350695469058,-0.00494864633580172,-0.0295041174501247,-0.0272880294777116
"354",0.0024996282136871,0.00200215008755067,0.0134730833090337,0.0034491397217804,0.00657905742228659,0.00333269653371304,-0.00401647398110505,0.00202615233162007,0.0108657378137615,0.00670297976193712
"355",-0.0103308615312122,-0.0148943041144282,0.00221567322820304,-0.0118970544050587,0.00385711019882584,0.00594187744117836,-0.0139685502894088,-0.0084556170451231,0.00583192701538926,0.0133169815653049
"356",-0.00583155867712093,-0.00295026751254479,-0.000736895308275143,-0.0180602543714575,0.00719840926839921,0.00525616848984378,0.000729642001291442,-0.0142751634124448,-0.0122783311991624,-0.023606741866913
"357",-0.000507070406454591,-0.00989345211095416,0.0117993756316535,-0.00871917640646735,-0.00890670561496221,-0.00363638309753711,0.00554641934904443,0.00921549800439347,-0.00264727219085892,-0.0149551263085738
"358",0.0199972850336987,0.0193312140269686,0.00801762356956459,0.0318167681241177,-0.00598962120665847,-0.00524799485508676,0.0251086335593751,0.00913181411028319,-0.0023081938301629,0.0379554310072467
"359",-0.0318938337647248,-0.0281265852873582,-0.0354305974891655,-0.0362303726638062,0.012946033290077,0.00871534641150973,-0.0396429920387723,-0.0232690882711617,0.0301908743848771,0.0255972879346751
"360",0.00242132796422534,-0.00103686674217385,0.00149947264654515,-0.00255703091743131,0,-0.00716268186047575,-0.0231461654497903,-0.0138019978068858,-0.0120143726030624,0.0102211742407385
"361",-0.00497737059772618,-0.0136831399336163,-0.0217065476377354,-0.0230703521072846,-0.00650041167515358,-0.00595522219225675,0.00392381956075782,-0.0279908342270972,-0.0277303677174762,-0.00400007566573857
"362",-0.0147123572506895,-0.0154994560585876,-0.0145371121025245,-0.014963701614225,-0.00232914779596716,0.00103813957003251,-0.0205955879534875,-0.00394469377620965,0.017182863219771,0.0368531702795376
"363",0.00380785601269928,-0.000874345661877496,-0.00232904526387512,0.00583171580953179,-0.0100039787102567,-0.0087463622967513,0.00614035740396424,-0.0128712841492932,-0.0163180768668609,-0.000227787839221172
"364",0.0126439356442354,0.00787889120451113,0.0101165599718052,0.0108080954858287,-0.00213367668529663,-0.00232097627391714,0.0208995039075939,0.00902712068321421,0.00268696267960178,-0.00638108513231939
"365",0.000587650921654248,0.00550056603263394,0.00924503560365464,0.00339913146498971,0.000224129998927181,0.000115533124656508,0.0143457859473286,0.00695827212737221,0.0137481064022347,-0.000917259715971785
"366",-0.00484456287762347,0.0012476362156506,0.006870232102411,0.00423401061545126,0.00202523099479412,0.00337381767845923,-0.0294642443660043,0.0059230518251272,0.0027582805939943,0.0101008964033154
"367",-0.00973665288150771,-0.0107362322898492,-0.0106140936308438,-0.00484892860850827,0.00842057520251016,0.00545083353975007,-0.014875150465787,-0.0107948380468479,0.0118051461318052,0.0136363564003168
"368",0.00126617594513023,-0.00164721018015634,-0.00306496330652828,0.00155371627741197,-0.00590049817596949,-0.00576680278180297,0.0206468967487168,-0.00297617752671087,0.00158585185303406,-0.0233182687419895
"369",-0.0162315540321769,-0.0198000887288361,-0.033051837580634,-0.0326447958511973,0.00582362370278244,0.00463982394170248,-0.024758059747095,-0.0107125422964754,0.00599410780353082,0.00688701191158803
"370",-0.000988288431438167,-0.00372095524310823,0.00715421746027078,0.00291539529866625,0.00211597081455017,-0.000461596731002656,-0.0207430801047074,-0.0207616381178229,-0.0209106358935571,0.00706784901461277
"371",-0.00197793106978972,-0.00377550485477429,-0.00789237622450323,-0.00443302921618249,0.00666607889772042,0.00531360210668552,0.000473907652922323,-0.0022861444880935,0.00436335994320181,0.000226438523680317
"372",0.00472612509932135,0.0134182353570089,0.0151877110943051,0.0200238963215336,0.00044161973080703,-0.000114435721257578,0.0176525636064329,0.0177083731046603,-0.000571658847928758,-0.00384796818793998
"373",-0.0271601779315691,-0.0245603367888673,-0.0251969412208602,-0.0343104604194363,0.0067299671113692,0.00563065387421702,-0.035759270804975,-0.0227222789504421,0.0364905407570473,0.0331744203459301
"374",-0.00545894288855198,0.00466271682681274,0.00565417844155558,0.00966901005454113,0.0117260370381111,0.00491370972789262,-0.00780686170934519,-0.00691289796352346,0.00949122602923258,0.00263902291314744
"375",0.00352840215321581,0.00268130985369774,0.0016066413664575,0.0075728712858012,0.000216464406562977,0.00068182528481997,-0.00327865213651801,-0.0101246844193797,-0.000765267292388017,-0.0177670229074153
"376",0.00312545730110569,-0.00874292950025712,0.00400957048697181,-0.017831006226583,-0.00236962026504217,-0.00271316352110107,0.00575648827374686,-0.0100145959179797,0.0137855795670552,0.0176417854465454
"377",-0.0171367289118545,-0.015357335668614,-0.0215655204209058,-0.0285068422550631,0.00522919180686299,0.00240020234503158,-0.0207685573749069,-0.00796376137081034,0.00550392810257172,0.0190915051542797
"378",0.00103043204317688,0.00779837165568886,0.00326535179180265,-0.00285753221355767,-0.00216680315372042,0.00034274372872356,-0.00801629394684189,-0.00282067643602513,-0.0119137063843235,-0.000430672741844051
"379",-0.0102129988310858,-0.0119209909872272,0,-0.00356223885748652,0.00456212628425545,0.00467445850293879,-0.0205387157945348,-0.000217286580772913,-0.00901580510570943,-0.013571687391414
"380",0.0177572043124472,0.00910147109884596,-0.00406812395270506,0.0122794598892824,0.00648695123056409,0.00249663900746344,0.0723615468477108,-0.00217644104041703,-0.00405570522671139,-0.0362524577358925
"381",-0.0192550059320212,-0.00985841907785334,-0.0163400688547592,-0.0201917990952445,0.00440412666268641,0.00475405408801222,-0.0735695980166152,-0.0071975688447784,0.00704379257050647,-0.000679765429519197
"382",0.00408690073383489,0.00646121536363364,0.00913612776745265,0.0181009129705274,-0.000107856441163068,0.000338112844382232,0.0181664560783614,0.00395435182091552,0.0221857814207651,0.0272107961405996
"383",-0.0116524099654284,-0.0181014693275593,-0.0131687109344015,-0.00669624794779611,-0.0142256909981525,-0.00934778481330256,0.000339760970264003,-0.0205692216998743,0.0174276169937733,0.0139072576091852
"384",-0.00904369699940866,-0.00321542593869406,0.00667222000372059,-0.0012396896267165,0.00878972302527026,0.0053428594589493,-0.0348221382493337,-0.00379766147334792,0.00788146246820243,0.000435523166912199
"385",-0.0140972388351387,-0.0148387082721269,-0.0165698420931774,-0.0166798209970431,-0.000322893753628706,0.00361884380087196,-0.00950390166219972,-0.0222020955784215,0.00271081210673296,-0.0317736170793276
"386",0.0245476995541112,0.0128792369208048,0.0252734658336937,0.028875990562206,-0.018076630580192,-0.00912615483360335,0.0701848184361789,0.0155959690882563,-0.0179889366328155,-0.015284340931413
"387",0.0100031020447278,0.0223062152833959,-0.00493012718655683,0.00467730756450924,-0.00514975676781293,-0.00477648652257234,0.0161045917080775,0.0219064298571692,-0.00232953192864194,-0.0235107378302527
"388",0.00623041637760413,0.00980263063852416,-0.00412879067245309,-0.00862447775960651,-0.00374523692990292,-0.00342790315426877,0.000326899478832576,0.00773460700861728,-0.000530704727969455,-0.0170640232062798
"389",0.000555515435951781,0.00584585172897589,0,0.0123954266068698,0.00387046452701623,0.00229316969869875,0.00294026289996308,0.0164469948491801,0.0100881917826949,0.0121285500252375
"390",0.0113447005789697,-0.000104032210217819,0.013267459255667,0.000608010072664422,-0.00495648175118513,-0.00343159814729588,0.0317591116456952,0.00539380046818394,-0.0216569063817208,-0.0218516034181685
"391",0.00541249570161906,0.00352893647607755,0.00654636549939802,0.00144407686223769,-0.00199288324238289,-0.00160717898296037,0.021309920682004,0.0313308287458345,-0.0267569100957857,-0.0225799169704837
"392",-0.0207537417596385,-0.0212016744894962,-0.000813031652907581,-0.0369584911084186,0.009759374604833,0.00862260631472211,-0.0615145938909772,-0.00728269315382857,0.00839132162967871,0.000737439518115224
"393",-0.000238853596972066,0.00612833729991769,-0.0113914361617979,0.00685556738653337,-0.00999416013506638,-0.00581325416660816,0.0151513768607396,-0.0253613688639336,0.00394174961257554,-0.0125246920014604
"394",-0.014663859220077,-0.0149128282375967,-0.0115227950903365,-0.0169050685350693,0.0100950516983112,0.00573298470229733,-0.0212524409947561,-0.0109678057143942,0.000436263487048283,0.00497402307860817
"395",0.0213521850997793,0.0110874892033701,0.00582884639947867,0.0554093889836158,-0.00406282800114643,-0.00284991954076208,0.0500583336756955,0.00217438312042773,-0.0124278530765991,-0.0113834159100783
"396",0.0178179009541448,0.00991134202375621,0.00910562598235742,-0.0104094701863132,0.000992079151114211,0.00194327427699936,-0.00489359909168974,0.0197439101000132,-0.0118114477011346,0.0197747231077408
"397",-0.0132265317235183,-0.0110669628345497,-0.0155863847070056,-0.0224103155585547,0.00991541746162516,0.0079874484478597,-0.011738732748339,-0.00531912268735957,0.00625564140713708,-0.00834558517007378
"398",-0.00528283368169458,-0.013091238983021,-0.0141665766963927,-0.00678376046675078,0.00221123565402914,0.000499671993725803,0.00240778254325358,-0.00342230953150502,-0.00566165617980341,-0.0111386394825681
"399",-0.00927393354931649,-0.00363737086224336,-0.0253592271586777,-0.0306166557357118,-0.00229362013051615,-0.00068148754418651,-0.0140911206240566,-0.0223226676570841,-0.0159651780730155,-0.0330412197272842
"400",0.0269623409545756,0.0300623911798867,0.0225498955672205,0.0128764643056065,-0.00744569030270859,-0.00511258249877178,0.0427155595676294,0.0208564519373717,-0.0233718745560686,-0.00698947251736459
"401",0.00444033418785073,0.00145922019301037,-0.00593722783683248,0.019909105669907,-0.00408226784667098,0.00034254835000036,-0.00467292165811217,0.00559108004514886,0.00650554120572644,-0.0106882484373897
"402",-0.0148915083724791,-0.0185263148524168,-0.0221842992481058,-0.0343371034935692,0.0162834046811433,0.00936060186643672,-0.0242567153788594,-0.0248073171801669,-0.00634814180918908,0.00553359520466379
"403",0.0185811529362554,0.000424413835264259,0.0148340046112698,0.00243565677023416,0.00272390289673141,-0.000452172169939535,0.0323977405587776,0.00197356100312174,-0.0192821010236776,-0.0280398631922217
"404",0.0103579203070234,-0.00190784419451351,0.00601878141993506,-0.0104472810479204,-0.00956450087381366,-0.0048651679095183,0.0245454557320479,0.00656614775873354,-0.0390856686012081,-0.00107836893611957
"405",-0.0104042477567942,-0.00488557886218177,-0.00683767787493084,-0.00834759934866391,0.00932825047589092,0.00693566167500226,-0.0221376733470464,-0.00478342791100028,-0.00751879727050897,-0.00863694178083629
"406",-0.00603059745599899,-0.0175027824351039,-0.0172114575644197,-0.000247602862745722,-0.00347920959016079,-0.00214499288569958,-0.0161267046322905,-0.0190081938859701,0.0129160586034298,0.0334875668411299
"407",0.00754435468213677,-0.00695175527801906,-0.00612948555996273,0.0131250378865178,0.00643694635794678,0.00305536592908662,0.0165486916989033,-0.0144767862314483,-0.0270966166526879,-0.00869334665424149
"408",0.00486334299676128,-0.00700066669352362,-0.00704876746058025,-0.0156437982757692,0.00867377110187229,0.00372244075991635,-0.00155047067108149,-0.00339001998155264,-0.0216761316112446,-0.0135530788405448
"409",-0.0136743132039751,-0.00638938226601327,0.00887345331524769,-0.0168857787720098,0.00397649008092316,0.00247306356581611,-0.020962653619083,-0.00680275774566796,0.0150715708516644,0.00565732592459312
"410",-0.010904361053494,-0.0121949587640928,-0.0158312478138131,-0.00833590629245962,-0.00385395846904169,-0.00145805726841719,-0.0206187133662493,-0.022830899205569,0.0206852403292421,0.0155371930081818
"411",0.00464605324895939,0.00224490547322698,0.010723902753645,0.0254714332614916,0.00279454803432788,0.00292026935245793,0.0024293065183163,0.0163548562420035,-0.00460029839612097,0.00791332262534139
"412",0.00172429875511937,0.00515096446918339,0.00618888754352098,-0.00149003563515548,-0.00182220814393841,-0.00212707849328952,-0.0137319871377782,-0.0114940690173827,0.0279790788903094,0.0429208050077479
"413",0.014475812476801,0.00713019897673517,-0.00702966029167174,-0.00074672994406666,-0.000643899783619339,-0.00291729496985826,0.0229319587502266,0.0090699840997075,-0.0148238269201523,-0.0338770128588113
"414",-0.0202853793670249,-0.016371873923633,-0.00884938912388411,-0.0206621075101745,0.00999136880711449,0.00663797171235503,-0.0220976978878248,0.00230476338944063,-0.00185004928835575,-0.00571443886543999
"415",0.00291283443471602,0.00382387204602463,0.00535692202382987,0.00177973885539418,0.000850938834215054,0.000336207245694276,0.00769626795573397,-0.00436903780015252,0.00370694427282814,0.000522586882356402
"416",0.00973421828488563,0.0109791295106587,0.00444065309947428,0.0213139927026871,0.00170041566902612,0.00145294886774106,0.0089374410371228,0.00808315431284412,0.00160036926257412,0.00939941240979691
"417",0.012127651445206,0.0141845439877004,0.0079571525073765,0.00695658502181407,0.000106160309212289,-0.00145084087014147,0.0331772498070351,0.0119128788959373,0.0100786503186008,-0.0196584834087645
"418",-0.0107535198894457,-0.00611898968346025,0.000877324077001695,-0.0118431951460081,-0.00445602324207683,-0.00122916984515131,-0.011223926375887,0.00271689388150098,-0.00571916524701888,-0.00369406808285622
"419",-0.0062117590875872,-0.0127529203571466,-0.0131462464845543,-0.0302120728212184,0.00930473705120649,0.00544340251363962,0.0122971966444916,-0.00541872134744847,-0.0307184191741331,-0.0259532462648115
"420",-0.00085918847855726,-0.00467697943394185,0.00444065309947428,-0.0164777676458648,0.00423936090302668,0.00245686891683095,0.0137049844547033,-0.00726415251906398,-0.00391411630987804,-0.00570970809837212
"421",-0.0301064959386026,-0.0449765390571768,-0.031830468761617,-0.0460733661184207,0.00801917325975188,0.0050113989753362,-0.0311872542952485,-0.0420767732902226,-0.00633793898260793,-0.0142191914588167
"422",0.00314471742490752,-0.00562320196070454,0,0.0142699915289932,-0.000523843002220303,-0.0022164531088551,0.00634306989270805,0.00501289246032521,0.00752652133596787,-0.00998620532375682
"423",0.0206554585981429,0.0172008771741994,0.0246577594428641,0.0124460117889942,0.00418939703049959,0.000111057200711473,0.0431770976047299,0.0261290101020812,-0.00151939725806294,-0.00224151519185878
"424",-0.0296876071088942,-0.0277971033402328,-0.0276293905549236,-0.056119898025603,0.00990866097554743,0.00455340667829685,-0.0438068402342127,-0.019907744651623,-0.0300532966008965,-0.0365066424621719
"425",0.00405831522671241,0.00428871248294138,0.0128324446561443,0.0161382924211084,-0.00619594132511647,-0.00254312096612808,0.00537090829266296,0.0243263839385699,-0.0296770435266582,0.00145725716199618
"426",0.0144678458935554,0.00142334361628205,-0.00542974949048536,-0.014767321253086,-0.000520486299740108,-0.00177307226152124,0.0114709557403336,-0.00806971546839463,-0.0153597276292141,-0.00844003600158705
"427",0.00462088945054107,0.0234544059271871,0.00636941891916298,0.0333708636673198,-0.0128922693022236,-0.00499614213122412,0.0105639134131399,0.016736196249614,0.0337985896606847,0.00675078805886775
"428",-0.0475848539872621,-0.0467593354223661,-0.028028898843431,-0.0785440887403678,0.0324418357168608,0.0191924257507003,-0.0614910923728537,-0.0477821772710875,0.026604830181145,-0.0393584528508193
"429",0.0167377508858384,-0.0118991489022418,-0.00930256531601337,0.00861295377684623,-0.000204852852473181,-0.00284694934714869,0.0307944134191764,-0.0177672504838569,-0.00992775941020507,-0.020333922337049
"430",-0.0449634377056746,-0.045956821531111,-0.0356806867531775,-0.0709656663581808,0.00500057588910074,0.00900361297757635,-0.0465596773116839,-0.0381325586661631,0.11290529869898,0.0300495994542949
"431",0.0296715505588345,0.0569291114278545,0.044790691650513,0.0843105905407147,-0.0146204691233788,-0.0117518891836952,0.0845001601345254,0.0200763214246358,-0.0311256263880836,0.0018046140202741
"432",0.039713747518811,0.0714108626885557,0.0540540495153572,0.124525141411412,-0.0317369302922433,-0.0178375801458949,0.0327338918550051,0.0652991799825546,0.0384057957099349,0.0330228692629901
"433",-0.0226393222043387,-0.02047301328105,-0.0344826139508997,-0.0652458467083256,-0.000106210895113645,-0.00212939927777012,-0.0880951660779349,-0.0179794915651653,0.0372179214741364,0.0345829335306627
"434",-0.0227515435991523,-0.0234552950217517,-0.00915796510052336,-0.0311455414726306,-0.00383205505645479,0,0.00636405432397091,-0.0158997590815263,-0.00964341780668332,-0.00983125370641769
"435",0.00320573053608442,-0.00190264994680089,0.0138634271540574,0.0114812158670423,0.00438145623654673,0.00258342987919558,-0.00739041022243359,-0.0061200196805612,-0.0182291779891304,-0.00822696864585204
"436",0.0156391456008349,0.0243029610423737,0.0173200828746365,0.051361710393625,-0.00202152559173541,-0.00302655388891182,0.0185310107066483,0.0187188546572503,-0.00299852384959665,0.0174484640515546
"437",0.000496895588057322,-0.00930442167165191,-0.00537652638102559,-0.0340080471130192,0.0072478451751159,-0.000673341984217202,0.0207925461108169,0.00580260642246544,0.00219782540883151,-0.0118076703580804
"438",-0.0783619623973812,-0.103545580552664,-0.0774774041102719,-0.116792218785436,0.0291001502853587,0.013946376213942,-0.0598346217425836,-0.0973556740488968,0.0338181098086114,-0.0620198269049511
"439",0.0413899793055337,0.0440025160970077,0.0410156415542433,0.0809867363154271,-0.0243697188714608,-0.0131998400008831,0.0485782010677334,0.0162452416459613,-0.0502400357262476,0.0279040396033075
"440",0.000603548749529725,-0.00125489258822475,-0.0121953064462307,0.011999126103444,0.0125805853184917,0.00704967559917602,-0.0153344820127987,0.00943396737469704,0.0105795345009991,-0.0233106248146986
"441",-0.0362743467963057,-0.0419492621312614,-0.0427348635694603,-0.0876230412326523,0.00803944235626441,0.00560046799986891,-0.0662297994436897,-0.0501039720428075,-0.0423403391608662,-0.0552870733393158
"442",-0.0135002304085911,0.00209777872987749,-0.0198413087382803,-0.0263073843568067,0.0088035636670849,0.00378675751524415,-0.0533706701591846,-0.0213173484036411,0.00315794963784888,-0.023345023034933
"443",-0.0509334309338147,-0.0580848254138944,-0.0323886010824155,-0.0751952906139518,0.0181726596957716,0.00810051369259535,-0.0183606925222485,-0.0823793590470423,0.0204625630445605,-0.0425672076916122
"444",-0.0447861664112384,-0.0500000664301598,-0.036610776729827,-0.0777897827809801,-0.00302529843782995,-0.000770455838052131,-0.0844508007942885,-0.00182568194565091,0.0354769581807897,0.0123118879564208
"445",-0.025192348766756,-0.0102340295612176,-0.0369163518871155,0,-0.0143620825918114,-0.012778698128776,-0.0167153935891942,-0.0423781388800176,0.0246361988530834,0.014527083835969
"446",-0.0698390277379912,-0.0747412056207259,-0.0462234727307558,-0.0736638589607006,-0.00841494807299703,-0.0100422589569488,-0.0715632299348244,-0.0799108074232855,0.00536797149111989,-0.0466200320130208
"447",-0.0242557638977985,-0.0249042994859816,-0.0437350761719814,0.0115369272216319,-0.00703630994523896,-0.0117223738526261,0.0795658951091078,-0.0311420192658212,-0.074304792562741,-0.0443590389076348
"448",0.145197813243679,0.137524656236034,0.158219997006472,0.227698445648615,-0.0128203154608786,-0.00684239300674294,0.0747487259681243,0.107142833172589,-0.0147801368086982,0.0555555194676047
"449",-0.014800245344366,-0.0184228360656959,-0.00533610937857576,-0.04976776000617,-0.00643956819863745,-0.00470846004554359,-0.0648741832044908,0.0438712336946885,0.00256127582781485,-0.0183518618979334
"450",-0.0984476067056942,-0.105571671603791,-0.104077325824267,-0.161661996368433,0.00956308815614459,0.00819128585925211,-0.141666771082328,-0.0908531130322574,0.0135036622933209,-0.0455026021484503
"451",0.0416571283570757,0.0498359307126894,0.0610777784091849,0.0491463003845827,-0.00515709006879894,0.000229913176714502,0.0628642945654154,0.0472468804421429,-0.0482534761314001,-0.0188469788539656
"452",-0.00597186355503576,-0.0162398209509261,-0.0135440042860739,-0.0313616605974704,-0.0068772297502977,0.00629216522801168,-0.0102766552761319,-0.032781621641272,-0.0262328411371821,0.0112994087772322
"453",0.0600795033025092,0.0520634726687559,0.0789475275682674,0.0700818275274318,0.00799045864616099,0.00102360114877986,0.00946018335981713,0.0620805777553837,0.0167076935203692,0.0201117479402557
"454",-0.0298554110094992,-0.0585395313191984,-0.0360551962160827,-0.0796631243989907,0.00528372499344387,0.0105629526022915,-0.0345142248625349,-0.0423379981160998,-0.0314649808917197,-0.0357795082209367
"455",-0.0544544176413906,-0.0762821322098519,-0.0605061147916494,-0.105284992279647,0.0202907606222467,0.00764283670414279,-0.0733900665194801,-0.0514679686673634,-0.0568196771908416,-0.0473305935845669
"456",0.0115843518376628,0.0183900955359495,0.0339579502725404,0.0279071627819261,0.00741884002836035,0.00133888776644153,-0.0155853508234444,-0.0285218681796858,-0.0147817182370898,0.00397460927152582
"457",-0.050714475460753,-0.0494037030429747,-0.0600226146588918,-0.103167699046605,-0.0106377888045074,-0.00423300601017274,-0.0641057687072408,-0.074829811134515,0.022080636317604,-0.0399841171555951
"458",-0.0355010169035509,-0.0580644979122779,-0.0602411090229161,-0.0262359274257586,0.000724152203478878,-0.000558749053752527,-0.0521350828666465,-0.0170280330983956,-0.000415441080396484,-0.00742275787031688
"459",0.116855544775861,0.129756407405619,0.12179501469768,0.209326374468313,-0.0145665125688913,-0.00805890036471402,0.163253290911058,0.0362204621876345,0.0223053615960098,0.0274200670797233
"460",-0.00725257315014471,0.0148197449463972,-0.0228572534722251,-0.0317052614484162,-0.00503154324158606,0.0014657783140315,-0.0397387790214324,0.0136777488303124,0.00284590048995925,0.059037684233568
"461",0.03459415121401,0.0288751588378855,0.0538011128977984,0.134956226106578,-0.00906120257582177,-0.00766143071047387,0.0484549662735507,0.0468516929373373,-0.017432445945946,-0.0412371829495353
"462",0.00550363990451919,0.0125803927063963,-0.00110991013524375,-0.00857742969687492,-0.0129720259771955,-0.00204364191592377,0.0629526630244464,0.0204080630244652,-0.0188420164879936,0.0111509323669647
"463",0.0028910199757286,-0.00382289084457454,0.00666662684671815,-0.00904420231376379,0.00270337231184836,0.00159847849243544,-0.0364277298770418,0.0245612517328011,-0.00336414372661309,-0.0110279603272104
"464",0.0339820652556382,0.0697155567244283,0.0551877856336327,0.0912697328553296,0.0187686784836505,0.0119713827587806,0.0556097746985142,0.0352740090137982,0.0616034475837819,0.0454003257497158
"465",-0.0420272854198893,-0.0594918678766143,-0.0209206682314618,-0.12727269115983,0.0118578072691276,0.00529582341984103,-0.0965803021030974,-0.0370490142945045,-0.0355060929184117,-0.0259048539988933
"466",-0.0554112841089128,-0.0632549829067478,-0.0865383196228724,-0.0504167558267562,-0.00721974986877671,-0.00302642460184954,-0.0452689142183763,-0.0398491420632702,-0.00796706011124759,-0.0438013163797875
"467",0.0330177038917667,0.0563285900453008,0.0584796812905737,0.0811759562980416,-0.00653400327839848,-0.00359791081054073,0.0592023244702717,0.0296962832294434,0.00387702847027116,0.00122699958366002
"468",-0.0131041650321967,-0.0215225576736183,0.00883963570798674,0.00933438012124377,0.00487953568771293,0.00101541186612497,-0.0857361283666905,-0.0535095858028658,0.0148965793103448,0.00653592119552315
"469",-0.030875572033642,-0.0252792140786825,-0.0416209199757402,-0.062323983893002,0.00295602448983967,0.00371936104595827,-0.0127251514160318,-0.0326726457399102,-0.0207936797827213,-0.0190745666179768
"470",-0.0440016222285399,-0.0565846788451937,-0.0274286767090256,-0.0741851130280218,0.00642120844734761,0.00617612988200866,-0.0736899169760266,-0.0288422491033355,-0.0284525040200208,-0.0293754072624588
"471",0.062339852059786,0.0828275129396723,0.0681551806375833,0.138489720477353,-0.0239525443180414,-0.00725365920929144,0.110708115943708,0.0441577407536358,0.0307143142857143,0.0187553871036426
"472",-0.0499069331485825,-0.0524233593732462,-0.0539051978339044,-0.0960128352126198,0.0198253114931777,0.00989124776207495,-0.0985838007120011,-0.0550149571358651,0.0159390293571995,-0.00627609242624128
"473",-0.013276290746263,-0.0327068421421542,-0.00232582275416837,-0.0166515374284436,0.00441307815264125,0.00422988104669719,-0.00785497912811028,-0.0213863748037189,-0.0088676804010499,-0.0227369028419511
"474",0.0188369889414748,0.0143883829064757,0,-0.0146453125163503,0.012867691770339,0.00775939841302775,-0.0401950152303122,-0.0129501490220081,-0.00192704743490579,-0.0150796573222827
"475",-0.0640790018128871,-0.0606381305984661,-0.0641026345555075,-0.0863913876468111,0.0256150345993287,0.0107790461976935,-0.120558478080523,-0.0873307608126732,-0.00344780020830782,-0.0113736460813515
"476",-0.0742325899193458,-0.0683277717170022,-0.0286425613635201,-0.0716825430733999,0.0516615751957383,0.0201302168628663,-0.0873017882736652,-0.0336926878971127,0.016468239234203,-0.050884855047417
"477",0.0539420515087623,0.0571312878026542,0.06153835906308,0.144030280645251,-0.0144600182501297,-0.00917310999494414,0.0826087778991256,0.0418410297728224,0.0735194175705685,0.0172494312916369
"478",0.0692914542734608,0.0770407414171292,0.0471015499385763,0.0607947693653297,-0.0156435267053852,-0.00936610073153998,0.144578433952437,0.0441769843349,0.0261256316074987,0.0687441540990277
"479",0.00740878831396174,0.0202850789638482,-0.00461374391067959,-0.0189530970977361,0.0294154976924486,0.0171701671420659,0.0271133566200339,0.0209401865904424,-0.000494388802650403,-0.0334477063449429
"480",0.0386415208042707,0.0177885206549762,0.0185401688462636,0.076357410575459,0.00134249827114186,0.00609009246468473,0.0456519061601302,0.0397657530492286,-0.00605918117747561,0.0319432230558587
"481",0.0125884226711106,0.00342697951998283,-0.014789517391351,-0.0192310928479835,0.0123522337509285,0.00201731919570647,-0.00861281461425656,0.0362312086460845,-0.000870850990452365,-0.0434221329352545
"482",-0.0885782715674428,-0.0877732754852889,-0.0577368645551929,-0.0962960888415745,0.0382954029617271,0.0135358995290686,-0.206111523985901,-0.0784767115566649,-0.0580251041719612,-0.0310112387636797
"483",0.0384848833214475,0.0490450752943785,0.0502449395488471,0.0631625326994416,0.00383950272377986,0.00524503062419757,0.137736073729869,0.0408934954025271,0.017184335302463,0.000463807880641598
"484",0.024041502352218,0.00749466893474793,0.00933502179619028,0.00816359120127208,0.0028224712067173,0.00156516661638006,0.045439472566779,-0.00648024229398969,-0.0100064591295564,-0.0115902577741106
"485",-0.0231332835322173,-0.0262129126797351,-0.0393061479411184,-0.0427352556716691,0.0197038318173288,0.00625211149506799,-0.0164975531990114,-0.0342439039263995,-0.00892622735626158,-0.052532722436711
"486",0.0308324928613735,0.01527811808072,0.0156436399985977,0.0592107949307461,-0.0162067759388841,-0.0105622010747494,0.0964515379183788,0.00253268947951391,-0.0129801721854305,-0.0247524516760373
"487",0.0349137423586561,0.0458618179222869,0.0450238653208814,0.0638860778518957,-0.00217197741519282,-0.00376752723214868,0.0941448367084046,0.0484209631763015,0.0225442843214285,0.0461928228227908
"488",-0.016483350450385,-0.00548143325269823,-0.00680274726266294,-0.0137613988815016,0.0197745395907394,0.0085091813163054,-0.0717927465531777,-0.000802953516470861,0.00170610242937408,-0.0218341123036047
"489",0.00681536754277223,0.0285910737315715,0.0216891303500444,0.0596194254945301,-0.00240073149975317,-0.000936518484233595,0.0663380124952238,0.0478294222442848,0.0448054226436416,0.0302580101527612
"490",-0.0240811256023193,-0.000669787504884778,-0.00335175138975974,-0.0255384687907962,0.00196150041073162,0.00604646466109449,-0.144254176155607,-0.00460301907014471,0.0112852915360502,0.0317765472120874
"491",0.01193947159394,0.00502670244152359,0.0224214017681394,0.0139231260509343,0,0.00279834942855839,0.094603263095191,0.00346864503342204,0.00198383132092173,0.0219319417556862
"492",-0.0139341729228908,-0.00200079329995517,-0.00548228679836626,-0.0133282865355361,0.0113908788720247,0.00217003650185132,-0.0284227210021692,0.0145923283863505,0.0221507244685244,-0.0282931297013179
"493",0.0470659446976092,0.0648182050198605,0.0507168280111758,0.0798200227428358,0.0247245345675502,0.0158814901248563,0.121791579813175,0.0264954184457307,0.0225181724580672,0.0143198584309669
"494",-0.00968675679321984,-0.00972714357631699,-0.00209879093809884,-0.0174373372552186,0.0271337969174563,0.00680173587499544,0.0252790094403401,-0.00921839407498237,0.0114847384736532,-0.0136472101417828
"495",-0.0186832264047776,-0.0323192488455438,-0.0347003424541275,-0.0219907620676691,0.0209827185225515,0.00675489637681626,-0.07889935986522,0.00446583343328832,-0.0182605290881425,-0.015267213431192
"496",-0.0043021610972912,-0.0216109358116564,-0.00435713048409592,0.00355023608360927,0.00106558961374481,-0.00330478445850402,0.0495912771754423,-0.00156733394754804,-0.0147848569887377,-0.00678285373721177
"497",-0.0128130447901899,-0.000576073234180963,-0.00218850979457197,-0.0373427066872677,-0.00768909090344783,-0.00261311282099086,-0.0209396324510598,-0.0332711320051288,0.0100448024946678,-0.0282925977976181
"498",-0.0103375773883493,-0.00576480657565559,-0.0171363077248726,-0.0082815737137395,-0.00131878646944528,-0.000503284462443299,-0.00759242972186369,0.0228152217572064,-0.0099449078593925,0.00401600906206068
"499",0.00580307869864716,0.0133013559389972,0.0123734019132649,0.00709816834233767,-0.00214576438683745,-0.0010080423040788,0.00765051572484055,-0.00189066074809296,0.0100448024946678,-0.0154999422095188
"500",0.00576993088670386,0.00807837550437251,0.0188889768460672,-0.00331662487821793,0.00330841322772635,0.00534739550854924,0.0132175501798593,-0.00378784827464762,0.0256410139664631,0.0157439728792961
"501",-0.00286836441142746,0.000333731522892844,0.00763355580142022,-0.00166403916327851,-0.00119931182931032,0.00220645071497771,-0.0563421703083925,0.0112020453065416,0.00876168244770281,0.0110000038080995
"502",0.0237027651977402,0.028371116031616,0.0281384433655503,0.0266664474590708,0.00952392544058189,0.00140728952904245,0.0452938413152952,0.011303466193346,-0.00521130295799199,0.00593463684071205
"503",0.0142745671840423,0.0107108726298064,0.00842108101380035,0.0133929667593877,-0.0209189324640289,-0.0110411917141919,0.0475523099437947,0.00894203367592628,0.00721763661891428,0.0417896661742048
"504",0.0301417771146999,0.0105970979289924,0.00521930962369654,0.0476571585314918,-0.0251361915147367,-0.0143102889694018,-0.0273971555350773,0.0347118997633888,-0.00335175693545164,0.0349221404623925
"505",-0.00118351129227978,-0.00953269834100368,-0.0249221681943944,0.0129968861791459,-0.0257840360328531,-0.00175016046892873,-0.0196081008853562,-0.00713805969231984,-0.0202945603515751,0.0104879131647666
"506",0.0066774977905304,0.0121912254820056,-0.00958510050571726,0.0226417027888552,-0.010057344156448,-0.00061941801711729,0.0495777468973706,0.0273186456404777,0.00769405749192509,0.0261732517063458
"507",-0.0299563943396356,-0.0117276266568577,-0.00967696705501819,-0.057564631112096,0.00392077378771893,0.000206876017308177,-0.0338167659573972,-0.0129459081921488,-0.0279572076103797,-0.0510114152463199
"508",0.00408102695946599,0.0128290300718974,0.0141151304244,-0.00430705309002799,-0.000798732721520423,0.0026829970510478,-0.00444435226605444,0,0.0206646404833837,0.0037070854943253
"509",-0.0214191502148889,-0.0345159147313906,-0.0171308039913455,-0.0216278783731019,0.00151063023993636,0.00463065290433584,-0.046037936740734,-0.0212692228247348,-0.00639357099684534,-0.0115419980752803
"510",-0.0240206449368513,-0.0272216311773992,-0.0119824577068351,-0.0422027997553172,0.0103783959528303,0.00624929561159115,-0.0582038329790632,-0.0315100627992356,-0.0376548626705163,-0.0453058901349086
"511",0.00184005345365335,-0.0188806430727988,-0.0187429987589545,0.00293757440194975,0.00105318338025495,0.000712427109192726,0.0301237968289922,-0.0373974055232711,0.00148582215240656,0.0166340748254159
"512",-0.0314545823325598,-0.0474229712737344,-0.029213626711862,-0.0485353209136814,0.0164887086952441,0.00559453455846715,-0.0518538287406153,-0.0470083779405369,-0.0134767067313318,-0.0139557828393829
"513",0.000356004521696818,0.00649363763934363,0.0127314981993796,0.0114333867319569,0.00163955064608245,-0.000809385438846122,0.0289346597323403,0.00163025441334042,0.00751971415566222,-0.000976072559683128
"514",0.00781985489686643,0.0014336596681257,0.00685738693227522,0.0108694847090567,-0.0154191699674048,-0.00921300326299901,0.0367737778297992,0.00488424264613174,0.0288593112185509,0.00439661793669699
"515",-0.0527867579432817,-0.0776664697728162,-0.0431330212158881,-0.0744086215690403,-0.000174770289046111,-0.00153239105999281,-0.108196323645697,-0.0810044837991033,0.0218836660849193,-0.0311282811770387
"516",0.0431926910370013,0.0364762755370478,0.0438911438324963,0.0543684427607871,-0.0315891773667138,-0.00890416976999009,0.0995986140993206,0.0599380592494367,-0.00437760308959789,0.00401600906206068
"517",-0.0154671672465957,-0.024335008932774,-0.0250002284631201,-0.033054727333845,-0.0192469954994918,-0.00660913045403766,-0.0507600226017005,0.0112268870615537,0.00510992263553356,-0.0129999764309525
"518",0.00435029544747079,-0.00652335388624437,-0.00233085376371234,0.0127620600759768,-0.00783049271881786,0.00020754121434341,0.0317004295708301,-0.014391289550728,0.0467013112626791,0.0466058108368732
"519",0.00685863325901415,0.026651245473311,-0.00116821925861665,0.0117014676118894,-0.00872929852562776,-0.00249342603864955,-0.00838015271708525,0.00709229497541219,0.004744131986266,0.00193618162824372
"520",0.0101580384329987,0.0161772767708959,0.0315787761217261,0.0177937071367347,0.0235130348105881,0.00656336460145224,0.0181537061335744,0.00289920992403703,-0.0064080946512004,-0.0270532163348416
"521",0.0338340363137213,0.0373935852287932,0.0181406155281416,0.0506994194776456,-0.0249861396463432,-0.00641739119535134,0.0796187666877797,0.0177617492305593,-0.0108621750688677,0.0238332003545942
"522",-0.0324981701247534,-0.0456815776461882,-0.0378619893120893,-0.0507488176234754,-0.0229978716555862,-0.0130224511510139,-0.0783031353887973,-0.0300329589403817,0.0237932057605399,-0.0121241352363949
"523",-0.020343071975002,-0.00710567735173007,-0.0243055247930273,-0.0074498191118928,-0.00317111239552359,-0.000422105974408948,-0.0318193370816467,-0.0121336906459981,0.020223441340782,-0.00589103658931234
"524",-0.00301841695990424,-0.0128057682545287,0,-0.0101546429267457,0.018605545149289,0.00811195777746709,0.00638126288730412,-0.00465909805040621,-0.0270507288807519,-0.0192592500730235
"525",0.0140474350396376,0.0335750123350051,0.0189800381224619,0.0298842576891964,-0.0238166780320378,-0.00861319946824057,-0.00380463816285259,0.0144682863569801,-0.00416473454141086,-0.0115811681446749
"526",-0.00489644306986348,-0.00996687366650839,0.00931307979201668,0.00736259793953797,-0.00349893064980777,-0.0050860065070788,-0.0235519199808307,-0.015100699048738,0.00802530792330391,0.00560380148302553
"527",0.0148810638995873,0.0193885996573422,-0.00346036464184596,0.0210660074660363,0.000877935908852878,0.0023426115330325,-0.0153192920643472,0.000425928213494409,0.0105405135680645,0.0222897741548633
"528",0.0284966458219491,0.0263350578528203,0.00578704777000749,0.0501052328453058,-0.0031186406120407,-0.00605626761483269,0.0685202449560229,0.0400169569623166,-0.00588112497066828,0.00743300010297254
"529",0.00137943783818284,0.00819669777487153,-0.0184119263258345,-0.00521241543404549,0.00322591620854262,-0.00203054273260139,0.0136310018396752,0.012280273811448,-0.0141756452361044,-0.00541064938474589
"530",-0.0458093456312465,-0.0516085325172126,-0.0351699818089071,-0.0604593446435894,0.021730805250771,0.0133886150412028,-0.0858803063707826,-0.047715490867745,0.0213994451992754,-0.0128586343260043
"531",0.00589580260586198,0.00782718261760618,0.00486042803947395,0.030029651126112,0.012971307237013,0.00771555015570935,0.0254097320528677,0.00127374930197943,0.0230573331455197,-0.00601204533501087
"532",0.000717890449481562,-0.00517763000793647,-0.00120936469438793,-0.00624695519560892,-0.00941548430501082,-0.00031441923081732,-0.0146725094054582,-0.00296877453632594,0.00953512829629299,0.00151228372584122
"533",-0.010758047462834,-0.0115239713187402,-0.0266344163556357,0.00502899046873662,-0.0266137124948055,-0.00786849103836085,-0.059894137811706,-0.0110585794143215,-0.00665444899977352,-0.018117878429032
"534",-0.0427736835543814,-0.0590450852134708,-0.0335823219179268,-0.0638032380987205,0.031149112327604,0.0168147885086667,-0.0630060438220215,-0.0692476654491599,0.03133434798484,-0.0558688131967552
"535",-0.00239900012254279,-0.0043962328474294,0.0077222844901228,-0.00712673854055212,-0.00852298175548849,-0.00728070740138809,0.00413221112212003,-0.0189461810496208,0.0152960402921751,-0.00597174427432889
"536",-0.0107552470600817,0,-0.0140485491193485,-0.00942152963440124,-0.0170004093867379,-0.00555245837301688,-0.0385331835201808,-0.0254359667242261,-0.0117635636461226,0.0245768480119914
"537",-0.00972056995092729,-0.0124446482848205,-0.0129534301456042,-0.0253622244948566,0.00971595646261636,0.0028441368879133,0.0642023639511522,0,0.0211966802087298,-0.0111942597399849
"538",-0.0357795074906618,-0.0402440262627926,-0.0419947753809371,-0.0246282637695402,0.00923806597367749,0.000946082711897001,-0.0760514577400998,-0.0362493098660187,-0.0007157463993126,-0.00970331719433548
"539",0.0379103700019163,0.0427784520432497,0.0410960916220613,0.0547882152490462,-0.00104852184636672,-0.00377857857860553,0.0823113563814759,0.0275826056723247,-0.0306968168209306,0.0190527660614423
"540",-0.00787309547468529,-0.0288384452566705,-0.0263159132333515,-0.0171636522628028,-0.0115497109323134,-0.00906005860765724,-0.0252286613499516,-0.0278183906893038,-0.0166789923990607,0.0117521957846016
"541",-0.0162610672975875,-0.000836131914668914,-0.0121621122306897,-0.00873157875891872,-0.0105247279470516,-0.00255218193762796,-0.0423856037963312,0.0115464488284442,-0.000966226495625944,0.0211193055324381
"542",-0.0223483964903841,-0.00711606344545523,0.00820785947884461,-0.0157628558831904,-0.00575768250315789,-0.000852387222806117,-0.0152762288345849,0.0143918145717341,-0.0046206856785016,-0.0118925004637856
"543",-0.0450428619708704,-0.0619731621757258,-0.0352778894428293,-0.0607629919745299,0.0165554442242317,0.0100326743133607,-0.0700081011509723,-0.0631116458452778,-0.0183525537629025,-0.0502355994577631
"544",-0.00750717729400185,-0.00898868813990406,-0.00281317861535169,0.0140425446908465,-0.00668170814815816,-0.00127089697727134,0.0038495221396424,0.00574409659360398,-0.0097877378203014,0.00661170746738571
"545",0.0236907595346019,0.0380953292982193,0.026798407196351,0.0702273879670319,-0.00458030902343698,-0.00508869540323076,0.0264172291942557,0.0150569592160876,-0.0116615169739948,0.0350300751350248
"546",-0.0408475458861879,-0.0397553826765709,-0.0192309336704583,-0.0411274412819459,0.0278101586502217,0.0117224869808719,-0.0643422358320148,-0.0424551075082974,0.033711653752369,-0.00846112494133433
"547",0.00174400071883052,-0.00136511510570436,-0.00280110911372899,0.0168673164164961,-0.00666943053351265,-0.00474031552248422,-0.0146407693851949,-0.0186964793587802,0.00326125672923716,0.0240000562089202
"548",-0.0117524905339901,-0.0241456763104482,-0.0351122170728579,-0.0194313211767954,-0.00585068998417415,0.000423544042213564,0.0211616584523229,-0.0446378995293576,-0.0186369160403412,-0.00572919525600046
"549",0.059609172960003,0.0732958877478145,0.0509461451735032,0.0811987469976443,-0.0191991034380375,-0.00729940779878691,0.132275266542244,0.0717947417825036,-0.0268300872253504,-0.00261919038814651
"550",0.00651267859700067,0.00521984670507147,0.00415506591646309,0,0.0108203283084745,0.00713958205589682,-0.0171341696176728,0.0159492427103598,0.012253256322365,-0.0315125524628562
"551",0.0393720424669801,0.0359151187798117,-0.00137934570413001,0.0384442983713824,0.00476797912144256,0.00285752286794794,0.0788429741573946,0.038723037467421,0.0210714747694298,0.0466376618266351
"552",0.00781441568154229,0.00167069034310696,0.00966855079029361,0.00559621715714553,-0.0050359423377645,-0.000738656071098021,-0.02129986501393,0.0292191200003977,0.00219544461460908,-0.00880838321565069
"553",-0.00302244198318724,0.0104253980193358,0.0177840282909425,0.000855917712214715,-0.0157696924805111,-0.00570183502850619,-0.073545911912609,0.0234947226767257,-0.00547645107963468,0.0219551233768189
"554",0.0305824282943112,0.0222865850372336,0.0349458852986433,0.0218135584711687,-0.00543948555059171,-0.00191196078722011,0.0745241692780312,0.0325205988127804,-0.00837006580275113,0.0214833462568833
"555",0.0223843739252645,0.0270487056843443,0.0233766849657724,0.0209291058666849,0.0378877893633951,0.0342624474943112,0.0516394650828806,0.0310330192697772,0.0338737779445382,0.0125188655265474
"556",-0.012386051537169,0.00353786180518112,-0.00507612160209581,-0.00655982134080479,0.00124551143566576,-0.00339503685431053,-0.0569894279397147,-0.00628963902275836,0.0135353104967368,0.0207713816451687
"557",-0.0212938707442628,-0.0117508629009405,-0.0216836233156422,-0.0136195381877996,-0.00555044467971932,0,-0.0744962934098092,-0.0134092817835234,-0.0080551353058852,0.0135659568000472
"558",0.0718288350924792,0.0729292343975132,0.0782270795442137,0.0924688277053707,-0.00866065196095789,-0.00340639032069578,0.149897649346226,0.0411019202154199,-0.0161341389522017,0.021032562538039
"559",-0.0197031358994606,-0.0369415577860798,-0.0278115703272275,-0.0310229650682626,0.0095134537471333,-0.00145031944679985,-0.071428619046217,0.00897257483605118,-0.0122719914797569,-0.0163857844833152
"560",0.0105460557420771,0.0149597767396972,0.0298508457947098,0.0150200948205002,-0.0134620939976462,-0.00601628551901778,0.0138825663064484,-0.00222276957039746,0.0113249701371623,-0.0152308792253397
"561",0.0203803970993284,0.0120937187204595,0.0108695194703741,0.0272584211765272,0.0115987855627386,0.0026085685979802,0.0248258360668352,0.016042751152358,-0.000543629032062398,0.0173997215694346
"562",-0.0180483066802481,-0.0403285846846951,-0.0167264053537252,-0.0295677927318129,0.00741842551690874,-0.000624440431701179,-0.0401208230987234,-0.00350866765312985,-0.0134885021211791,-0.0185273076455011
"563",-0.034554636220661,-0.0412452143025946,-0.0388823024085141,-0.0515623778272277,0.00382607390667555,0.00427009034928516,-0.0548108842198965,-0.0528171751198064,-0.0078288563716209,-0.0363020355662409
"564",0.00926508972484608,0.0381491494305963,-0.00126410449317971,0.0218285668709286,0.00714525758272466,0.00176361161793381,0.0621609999161008,0.0250928958669221,0.00333402967323759,0.00452038323437498
"565",0.0193662658213185,0.0234561216670568,0.0291138798100663,0.0330511104246944,0.00912616569121405,0.0024503636005182,-0.00903422124840758,0.0117860009229638,0.00830748790770364,-0.00249996577856626
"566",0.0292377515227238,0.0469822407967126,0.0356706146405892,0.0542334892952243,-0.0122210581201627,-0.00652486369559069,0.0661911966231246,0.0640684326174332,-0.024497374761039,0.0385963742912467
"567",0.0099486593289968,0.00839127941885498,-0.00831360943605863,0.0122129943998104,-0.0204621940467099,-0.0114683113086452,0.0895909992104877,0.00505228891011855,-0.0136262044946103,0.015444053609444
"568",-0.00783290579109508,-0.0188132953445668,-0.021557151427733,-0.0124313912747096,-0.00427577992792738,-0.00232043389191838,-0.0160352389525992,-0.0146627554763348,-0.0264870316925234,-0.0123573436304513
"569",-0.0233254136124222,-0.0265487954133601,-0.00611992672128725,-0.0229545750613867,0.00253760090948152,0.00253760957313554,-0.0752428519789082,-0.0153060990739696,0.0172393696694981,-0.0178056351805647
"570",0.0107773183857387,0.0102273739629903,0.00738946314561528,0.0147783901251968,0.00885672000553783,0.0049546455269176,0.0209972941860535,0.0250430514315267,-0.00149869729072394,0.00734928855250017
"571",0.0397427078228816,0.0217475506248983,0.0366745498140268,0.0436894162074914,-0.0125421626997323,-0.00587492799016376,0.119353854748603,0.0421233407865995,-0.00346383785401416,0.0145914913061271
"572",0.000233804248785274,0.0176143823753199,0.0023585512868296,0.00608219609791849,0.00918463870933905,0.00590964673920391,0.0127949414551511,0.00525459400476636,0.0181902333029831,0.00431451718146958
"573",-0.0172435805453562,-0.00937609290186214,-0.00941155091469736,-0.01600282524381,0.0052274918479378,0.00514153421233754,-0.0819564615014419,0.00723754995487647,-0.00580330015259334,-0.0181385200973956
"574",0.0106700772403923,0.0152894945315916,0.00475046720078898,0.0144561821960447,-0.00173360839578163,0.000940398744784465,0.0818632189625659,0.00518942199582617,0.00148789052920151,-0.00631979731497179
"575",0.0146621226081232,0.00609542462108448,0.00354576757420144,0.00854995568322581,-0.00791091704636826,-0.00396382603349343,0.0407694302258552,-0.00198530924830909,-0.0193143085714287,-0.00440312116309871
"576",0.00670560349630667,-0.0017821900213203,0.00471172276483567,-0.00706455400821548,-0.0109891079442956,-0.00806197686015309,0.0100283384381041,0.000795310957645068,-0.00687562071729675,-0.0073710074952722
"577",-0.0419153861595414,-0.0485539519269844,-0.0222744777781957,-0.0487371026005685,0.0151426726574693,0.00696677657086453,-0.107042988764475,-0.0588466182500491,0.0203003517918288,-0.0376237562217255
"578",0.0195374382034681,0.022889458873167,0.0119903954268781,0.0213161890920102,-0.00988056907291268,-0.00387862269860895,0.0913826717864108,0.0190116468337236,-0.000690028775964135,0.00360077366973188
"579",-0.00611318135646155,-0.0110051174468814,0.00355466464553267,-0.00842169254219738,-0.00606495368447035,-0.00242025869237938,-0.0337469275141302,-0.0037318286884368,0.00563929112256067,0.00153775748535745
"580",0.00981744164616027,0.031527879309436,0.00590333905164542,0.0155095288937293,-0.0000984579196280366,-0.000210508104872775,0.0415153603755845,0.0228882330542193,0.0162509275435201,0.0133059086425964
"581",0.0151107602940446,0.0172602443565735,0.0152581153945908,0.0189092036734326,-0.0100400185686441,-0.00390388543051767,0.0528313607484081,-0.00325450859037935,0.0103603374878263,0.0151515687072972
"582",-0.00946213323423273,-0.0130788639161648,-0.00231240448195202,-0.0335475042586449,0.00427518451367814,0.00413056310350268,-0.0564906275047659,-0.0191840099629855,-0.00791349745972469,-0.0248755890277783
"583",-0.0031454596583339,-0.00286536472722487,-0.0162225539471361,-0.00332354646937882,-0.0163370706450604,-0.00485246369234904,0.0108283933339719,-0.00457691696732798,-0.0141557349925686,-0.00714296929139702
"584",0.021269147895147,0.0312499111169418,0.00824545344450955,0.0526121525565391,-0.00885622185495671,-0.00540593167521641,0.0396973683983499,0.0292639680669251,0.00660970940170924,0.0231244135623185
"585",0.000343215753374704,0.0045280226289357,-0.00584140945128142,0.00915162871028774,-0.00396104261803099,-0.00170499501016674,0,0.0125913212589943,-0.0120005091814669,0.00351577321474195
"586",0.00537642498740221,0.0124827699287908,0.015276224224001,0.0146494357749045,-0.00688285526570032,-0.00321195148349018,-0.0339391329417044,-0.000401102104038875,-0.0036667813796305,0.0300301367672682
"587",0.0340194785014607,0.0410957307408155,0.0266205024776738,0.0690959964329105,0.00329544777975865,0.00096665064198187,0.0865743390157849,0.0389245681163635,0.0194364814066641,0.0194363296856011
"588",-0.00341086665500911,-0.0108552386407323,-0.0033821056791169,-0.00900324068815683,-0.00123218352817267,-0.000214568798088455,-0.0334871148054303,0.00231737546963884,-0.0043998082626332,-0.014299382269237
"589",0.0173344529816606,0.0216163824367239,0.0237555536567544,0.0171967540770037,-0.00236342268979584,0.000429229695476652,0.0334528628004063,0.0354531895955124,0.0146175750708215,0.0265957801542649
"590",-0.0138916734035704,-0.0179036625557577,-0.0232043221371565,-0.0248805670689352,-0.0244128389548528,-0.00836896283548816,-0.0578037551317296,-0.00744380425338298,-0.00111680811797177,0.00188410047824861
"591",0.0233324040800058,0.0477294759040441,0.0407237051890015,0.0333663143568907,0.00242918883909016,0.00118999172732126,0.0677919098125599,0.029246598565035,0.00603757812974992,0.024917674809716
"592",-0.0187132596543956,-0.03068640979632,-0.00978240723279322,-0.0234253236595574,0.0142193480711041,0.00940261538883025,-0.029301941745112,-0.0280513940997879,-0.0032229494368875,-0.0082568156770203
"593",-0.00295940596245337,0.00979110700055186,0.00548825470858527,0.00713150066080015,0.00363469982615316,-0.000643242451454307,-0.0159814106657178,0,0.0112609541473752,0.0101757669694855
"594",-0.0251729054697455,-0.0303816672903978,-0.0185590071999955,-0.0366915328363863,0.0108643680686644,0.00460750603067273,-0.0679699888225105,-0.0431028487013334,0.00429987886328154,-0.0114468713857856
"595",0.00857002387954098,0.0103337644779671,0.00111247515418045,0.0143669037776575,0.00389051192507583,0.000106248631053241,0.0319459645966378,0.00940042469777147,-0.000658656302937932,0.00648449018123598
"596",-0.00816206290354116,-0.0131971711200662,0.0100000913401466,-0.00922256306055913,-0.000305541486430916,-0.00245234717492715,-0.0328328150150168,-0.00388049055784856,0.00571244650897995,-0.0253106155559778
"597",0.028406985659418,0.0434636122510601,0.00880087594262102,0.0555184865414908,-0.0155039941169143,-0.00587918194458703,0.0750077450859219,0.0268799260280692,-0.0129983829711071,0.0264399184207804
"598",-0.00120541475723612,0.0124962176578027,-0.00654301534906043,0.0113384733286714,-0.00528361284173695,-0.00139777436855126,-0.01593950915215,0.0170711833967765,0.00664008403452754,0
"599",-0.00669457018284936,0.00474678376000748,0.0131722167142636,0.00311449030678368,0.0105186071439729,0.00312286354008751,-0.0116137354683599,0.0104437244256279,0.0141820691972523,0.0160994686754468
"600",-0.014363508042848,-0.00440950312921207,-0.0130009651833735,-0.0186279111288238,-0.0251488573345955,-0.0109494267366528,0.00185539115925204,-0.010335780383578,0.0173441517615176,-0.00814846504239086
"601",-0.00212940100422354,0.00379622607312946,0.00329313591519065,0.00442905025506635,-0.0111016684187132,-0.0058606072502625,-0.0212964971878633,0.00522213470637389,0.00319663299300221,0.0146050497443448
"602",0.0256120090439251,0.0211157722642228,0.0328223878122322,0.0119686076938175,-0.0150755619675154,-0.0066586205600081,0.0517184274704308,0.0330233940952309,-0.00414232598741737,0.00224927486095283
"603",-0.0178533279520944,-0.01697528171189,-0.0190676583039537,-0.0115157914262588,-0.0176944934882503,-0.0113205958474446,-0.033282856798536,-0.0114937861116107,-0.00330636725029088,0.0044882691767838
"604",0.0139401574400719,0.0128728032230729,-0.00647951950312986,0.0308563701483406,0.0144764665607169,0.00522501722348778,0.0189204693764038,0.0148976728218115,0.00845372953837553,0.0183200938637791
"605",0.0177080088869428,0.0136391773775599,0.0184783803396797,0.0152720318964594,0.025817655113954,0.0112791181021483,0.0273970756749962,0.0329402008269559,0.0207979524787341,0.0193066290542936
"606",0.0242078297535513,0.0284403987373192,0.0160085665871632,0.0421177389278784,-0.0295636400538726,-0.0163194030786156,0.0420743109801456,0.0183705504980118,-0.00488559266794986,0.027550648242207
"607",0.000844387108655642,0.00713632513334894,0.00105044705086721,-0.01443421796976,0.00537845791316327,0.00334490720474268,-0.0147853741796578,0.0139553986969483,0.00658098798973183,0.00418930158616559
"608",-0.0126511864586134,-0.0345437204093545,-0.022035646343403,-0.0354419973566668,0.00939112004589648,0.00611159861896726,-0.00230897504346261,-0.0184626423964909,-0.0202365813591056,-0.0333750258162775
"609",0.00939644271071893,0.00795091339598586,0.00751063377411998,0.0185238235093743,-0.0206620542751063,-0.0115967624621848,0.029505462827226,0.00273583438982561,0.0192776074874437,0.0366854001460537
"610",0.000211642550440372,-0.0127425823865505,-0.011714731630286,0.00208705681927501,-0.00762106207212587,-0.00994579168934462,-0.012644109080702,-0.0225099870489631,-0.0261873004410069,-0.00541225372086029
"611",-0.00412503445393775,-0.00522438238650458,0.0053880378011899,-0.0154715286863936,-0.00256096100185121,-0.00507901683194256,-0.00369965155023577,-0.000349282342996915,-0.00160069364636317,-0.00251151998290522
"612",0.00509805606226021,0.0120481488208191,0.00857455134963758,0.00181335794803106,-0.000111284985618743,0.00431030755090012,0.00114294245634072,0.0150088976677369,0.00288589146827478,0.00965169779847508
"613",-0.00253615160720122,0.00274722327328325,0.00106253655446698,0.0126696603467873,-0.0157371699883077,-0.00598623516106234,-0.019115703046789,0.00447063160813532,0.000319716501764544,-0.00374059749461575
"614",0.00444933189817553,0.01674299982856,0.0169852278927056,0.0214476988715422,0.011113151784397,0.00681827792691014,-0.0186155852335309,0.00581955575569459,-0.00170470912311205,0.00917814283389506
"615",0.00274181915689775,-0.00508986180252002,-0.0010440235960526,-0.0160396438540866,0.00897129451281109,0.00530544263831922,0.0281564443889777,0.00646714356253075,-0.0163286984950489,-0.0140553730163712
"616",-0.0229278631331216,-0.0373158020197218,-0.0177637445657457,-0.0358624668998199,0.00900260936215758,0.00449002850142688,-0.0449697087273737,-0.0246870619324114,-0.0116089836521425,-0.0192872499722414
"617",-0.0135628840587237,-0.0128162949378046,-0.0106386036084579,-0.0150631072587546,0.0174052586473115,0.00558918679743892,-0.0141863224192069,-0.0149099503316186,0.00911088933284065,-0.00384783372232922
"618",-0.00098201773736073,0.0031662917716444,0.0118284254746104,-0.0112358856509557,-0.00563036018674712,-0.0026678405666859,-0.014084221671632,0.00457593496643693,0.00456867181551179,0.00300442766130105
"619",0.00731786263482337,-0.00315629801122252,-0.00850165348527121,-0.00284084191850309,-0.0151354728118039,-0.0121480275906234,0.00496870025447516,-0.00455509116549735,-0.00801296173281996,0.00128359132876055
"620",0.00368624793507344,0.0145657867521098,0.0160770084384925,0.00506474301412507,0.0137102733947145,0.0046257438884747,0.0108155788486781,0.00997114100919094,0.00316560415712686,-0.0085468920092806
"621",-0.02998710330563,-0.0362211551102113,-0.0221519367148924,-0.0362204562871901,0.00970636485930343,0.0053897361898918,-0.0510548381921045,-0.027855824121545,-0.0147987047921936,-0.033620804004005
"622",0.000784169822614755,0.0201985666026792,0.00650774566384849,0.00649001903319735,0.0117731413973996,0.00323938350700304,0.00869874568668516,0.00652900597134676,0.00419700680144675,0.017395175235059
"623",0.00861780355558728,0.00194736672680018,0.00215499945380415,0.0219314007476987,-0.0100347635240579,-0.0037853372270138,0.0164379681416496,0.00504472764162722,0.00582928961349061,-0.000438398234711701
"624",0.0217487352432888,0.0129576231729216,0.023655930830268,0.0297887778793828,0.0183323834008973,0.0125168567072111,0.015949047177555,0.0340627060068148,0.00940405717017123,0.0087719456635289
"625",-0.00260652248455528,-0.00319775049099835,0.00315152154104514,0.00528769472818924,0.00169443373960365,0.001324968583585,0.00879117901017556,0.00970862787108784,-0.000216628755641324,-0.00826089106396555
"626",0.00936409845287622,0.0112286631818617,-0.00523563116541537,0.00742584477389086,0.0014802519244268,0.002094050532091,0.0024897765390226,0.00583774031450335,-0.00270885250071673,0.00964489652745826
"627",-0.00809033300387441,-0.00444187661495998,-0.00736840605180156,-0.0101352974459106,-0.00168916849468392,-0.00263994859200734,0.00651964666106486,-0.0191188804051676,-0.00934377434437439,-0.0178027572355389
"628",0.00413268177358317,0.0152965593370658,0.0116648887971855,0.0183057889121763,-0.0019844073277735,-0.000641563722688199,0.00987048495641063,0.0156631618154752,0.0132704430796227,-0.00397881616864659
"629",-0.0272935427592,-0.0310735590804828,-0.0220124094871148,-0.0274221657446063,0.00233902195120672,0.00331975554560549,-0.0455099199283777,-0.0215905023392395,-0.0123389870368978,-0.0221926019969989
"630",-0.000110909108948842,-0.00161957086279385,0.00643069971056254,-0.00219275487817117,-0.00190835507136022,0.000662179815823505,0.0208000597689362,0.00910673863503941,-0.00536984109589045,-0.0299592023076115
"631",-0.0193766410177373,-0.0295262188725663,-0.0106496550486995,-0.0235482738638931,0.00669365326021976,0.00396823936787394,-0.0369904749753599,-0.0357512180695353,-0.000550936523778467,-0.0159100812892855
"632",-0.000680835267292235,-0.00668689239904308,0,-0.0115753451365109,0.018469592639055,0.0115287002075184,-0.00976591768338364,-0.0104390756523675,-0.0158747879602555,-0.0123634141565601
"633",0.00193125714587361,0.0151465299264681,0,0.0178918143645745,-0.011917390078297,-0.0058620307595818,-0.0161078203508445,0.00800265082719509,0.00268852927148622,0.00625904125719567
"634",-0.00238190011528205,-0.0079578382104889,-0.0107642272585805,-0.0118247561630231,0.00922947288013254,0.00622370128251393,-0.00167082382414219,0.00360904481352242,0.000782035509282908,-0.00765554569948457
"635",0.0243291627313877,0.0257354245007075,0.00217636158954382,0.00711534484047971,-0.00561207089516413,-0.00358074154364862,0.0394914373348341,0.00898938719003239,0.00680955555236551,0.00530393685595221
"636",0.00566073512517251,0.00260693673246815,0,0.0109182326377255,-0.0166161800487485,-0.00664238227532343,0.0115902819179396,0.0242336535597498,0.00687433181340857,0
"637",0.0292460670525827,0.0425737946362419,0.0108576941507599,0.0536848967162606,-0.0257172717729671,-0.01293636611301,0.0343733654433567,0.0208768309184475,0.0157471647560217,0.0263786816745606
"638",-0.00160820107627546,0.0109101041048647,-0.00429661927371194,0.00180880414289875,0.0107987184893243,0.00599756846303912,0.0129232647352755,0.0248806379462705,-0.00281867959277282,0.00233656119252856
"639",0.0109544462113462,-0.00370017730033678,0,0.0102318322665111,-0.0154309778342433,-0.00673467772161573,-0.0233901823752054,-0.00897898524001517,-0.000543629032062398,0.014918402839005
"640",0.0106235152075262,0.0194985607416231,0.0129451280908695,0.0357464719013676,0.00526127908849827,0.00366811491326779,0.0323482655584966,0.0218124988793382,0.0146850756010006,0.0165364813130622
"641",0.00462528062137912,0.00455383732603187,0.00851980606543523,-0.0028763047449345,0.0199521380509344,0.0111852088971762,-0.0021092427553927,-0.00426921992268636,-0.00160808320763384,-0.00361499950632049
"642",-0.000209150491115473,0.00392852443117997,0.0116154290456298,-0.00230757387684022,-0.00897954279375535,-0.00591392541565194,0.000906136895489906,-0.00428776245636431,0.00332873413493195,0.00544224272584604
"643",0.0220828514674367,0.01745963868509,0.00417537044449379,0.0283317150367384,-0.0183370598066971,-0.00969488875003199,0.0346907069416131,0.0215300563765404,-0.00192636982178152,0.0207486147016711
"644",0.00409582724002377,0.00739624063692479,0.00519750382104189,-0.00477908294870544,0.00483479189276825,0.0021138805270926,0.00874622678290793,0.000648492905181097,0.00160842801611771,0.000883861571832734
"645",0.00295719231348457,0.00146843546066133,-0.00206827016296107,0.00875702076182061,-0.0114816216928896,-0.00466255124719805,0.0187862713686966,-0.0116653074241551,0.00321159391021975,0.00397354664689109
"646",-0.00467717426499847,-0.00586500975144277,-0.00103601744676962,-0.00448042575961749,0.00884947730049501,0.00200686879463041,-0.00397161796371504,0.00557348760206922,-0.0170739303924227,-0.0109938289580486
"647",-0.00245161625515378,-0.0097346287188681,0.00726130268981029,-0.0225034758653664,0.00548193513743556,0.000668548812277958,-0.0142411166306999,-0.00912928288098935,-0.00987953523092455,-0.0257892071251772
"648",0.010445249406938,0.0196604846461275,0.0113284252389072,0.0247480309442458,0.0141769674781087,0.0040044200763194,0.0349610433852947,0.0164529782275511,0.00460532909885947,0.0310360066831867
"649",0.00141898679191144,0.0169441898036939,0.00509164821993391,0.00477385344369718,0.0194621854080765,0.0100817888376337,0.000837583971234013,0.0213657944272918,0.018882284908897,0.0199203653748934
"650",0.0164963873740616,0.0264293138593281,0.0172239238866898,0.0374508745520838,-0.0151547830536427,-0.0106262446469463,0.0198046707276456,0.028843187951898,0.00557048753230815,0.0282116866853799
"651",0.00258829663335236,-0.003358734691292,-0.000996009735260595,-0.00915925261617978,-0.00795099456948523,-0.00289129564970103,0.0475930140681946,0.00462082203917991,0.0086289227028149,0.00042220018779604
"652",-0.00287996206077856,0.000842532528478213,-0.00697884210457611,-0.00842845488529287,-0.0149489719254137,-0.00568628767451862,0.0404699544803981,0.00276018380337528,0.0010561787072243,0.010548596042903
"653",-0.0051783275495465,-0.00841766083682871,-0.00100400958407387,-0.00822584043290242,0.00340942613162531,0,-0.00627340880306371,0.00152909799117285,-0.00189914540936009,-0.0229646233327346
"654",0.0131142458441116,0.000283105201185574,-0.00402010430268906,0.0099529480201539,-0.00832928821296175,-0.00661694101238808,0.0464646696284767,0.000915484806226496,-0.0089851798939784,-0.004700702637916
"655",-0.00207503512432761,-0.00735488546477925,0,-0.01122379436378,0.0124879315660111,0.006434637291858,-0.0197879863512874,-0.00274504376887397,-0.00874666666666657,-0.000429451290466343
"656",-0.0124761728234228,-0.0108292972653599,0,-0.0188261747615885,0.0115693536023964,0.00695480522132197,-0.0295418187033993,-0.0171307602790252,-0.00150649951576454,-0.0150343792638081
"657",0.0107286876027712,0.0146931426990529,0.00504540599344505,0.00902964729462052,-0.0106821069809852,-0.00278491331894548,0.00659554978678312,0.0289451447397695,0.00172428061510632,0.00523324715238638
"658",0.00763908048742268,0.0167518194310319,0.00903614574295442,0.0173374809428881,0.0141780786043626,0.00781993265826286,0.00478849067317788,0.0057469055145154,0.00828406696990003,0.013449063960312
"659",-0.00767978496543442,-0.00949457411986543,0.00397966113425685,-0.0181414847625702,0.00387178441063107,0.00310382855877434,-0.00902949724217295,0.00330838139755629,-0.00768246897479219,-0.0282533912361369
"660",-0.0246053363735754,-0.0352411298298992,-0.0277499633074083,-0.0391937958847243,0.0147830177620396,0.00685073128940639,-0.050113835516355,-0.0344723224840922,-0.0149462258064517,-0.0149779951796416
"661",0.00793398324835759,0.018702495166786,0.00815495286177526,0.0218531895441556,-0.0058057958090304,-0.00351257255490955,0.0122571971014025,0.0229740122840343,0.00491209469586185,0.0196779575566206
"662",0.00877996290923155,0.00975343707363829,0.0030332580048551,0.00256610531614521,0.008281540492594,0.00374441892470134,-0.00737068880165115,-0.0145673965339568,0.0051053770390046,0.00701749333334312
"663",0.0103039991760039,0.00909072557790225,0.0120967886434278,0.0173494001790182,0.0082141649549643,0.00263383258130467,0.0405726240194275,0.0163226162619066,-0.00280992113703582,-0.00827519375240693
"664",0.0196055636596326,0.0295609091486313,0.0109564316555593,0.0150965792376236,-0.0205766105898395,-0.0101774661708863,0.022171396798113,0.0148487581607533,0.0149561617521241,0.00746599767470402
"665",-0.0000967465393496569,-0.00136720994323969,-0.00197057651438914,0.0044062517205905,0.0181290018491076,0.00619081031857505,-0.00573431342015773,0.00507609999549929,-0.0139883179073504,0.00174365530253318
"666",0.00194245877077037,0.0076669099696951,0.00789725528947249,-0.00219337574632006,0.00565714155110131,0.00263758119583923,0.0110333162374079,0.00950644220591967,0.00454847323146956,-0.0143603410888363
"667",0.0000970976594085737,-0.0040758473325867,0.000979425791174604,-0.00302315284169741,0.00458191079487991,0.00131474580131963,0.00446417487951845,0.00176623377727259,0.000323404477718725,-0.00264897051125457
"668",0.00222897548072853,0.00818550054663914,0.00293554729711554,-0.00192930637062549,-0.00393929693878414,-0.00273539845931181,0.00790122428071771,0.00793157269195044,0.00431082008502193,0.00841077740029217
"669",-0.000193408542298656,-0.000812198367161066,-0.000975748032788659,-0.00524713495745999,0.00458056697013354,0.00230445824871395,0.00661468181608438,-0.00058306427160304,0.00729693084457694,-0.00219496822668053
"670",-0.00889893416368082,-0.00622963414666899,-0.00195311279521482,-0.019711247162584,0.000932006817067066,0.00295594994024428,-0.0124119430597516,-0.0067075190155258,-0.0050069349630254,-0.0272766279455596
"671",-0.0220576393419685,-0.0283454486624086,-0.0146772437155004,-0.0189748768219653,-0.00241991297917898,0.00259456362763721,-0.0510104134808554,-0.028478925706277,0.0053533189431838,-0.0153776794646028
"672",-0.00379242950112835,-0.00364668692197334,0.00297915716702213,0.0106815181779178,0.0145749972977953,0.00545996859443276,-0.0197353457471741,0.00604424928372693,0.0243876459129362,0.00229675452761691
"673",0.00831499095699595,0.00760150887277455,-0.00297030815220234,0.0199941264099499,-0.00615740565999712,-0.00358445745719571,0.017748305925805,0.0156202535571786,0.0132030041957998,-0.00504131910971206
"674",0.014009108579639,0.0192792294989355,-0.00198576156505115,0.0193223819237547,-0.0170342333224242,-0.00599372532331521,0.0119731445469813,0.0201124941816393,0.000718243389270068,-0.0041454986395717
"675",0.00862243567793053,0.0249449342365327,0.00895525450126033,0.0206044365379321,-0.00703740346636417,-0.00230293715499197,0.0321501052311473,0.017106594566507,-0.00102531529811656,0.0185013728514223
"676",0.00767435275004846,0.0117680663830251,0.00394465994519355,0.0053836708295063,-0.00116290413319098,0.000878962628548363,0.0201842774119578,0.0188140909083658,-0.00359230216565753,0.00408723115819432
"677",0.0102187693115487,0.0113665033643726,0.011787715029528,0.0131189773079219,0.0184262402130886,0.00746651264761211,0.0141672026916906,0.0125905516010782,0.00638643373740355,0.00542728758512201
"678",-0.000190653524230089,-0.00313627865835875,-0.00097109778975446,0.000528458234429374,0.00551101455823333,0.00294320173557994,-0.00313119676927598,-0.00442115426169643,0.0110542685072959,-0.0130453034291789
"679",0.00486783952275083,0.00498171819246385,-0.00388692900968801,-0.00369735225195167,-0.00992800931420812,-0.00586827919848343,0.0287512171335915,0.00471840265716783,-0.00830127564589267,-0.00546948107058731
"680",0.0041793579199727,0.00391315246559887,-0.00780511721331834,0.011929647817122,-0.00511720675493244,-0.00207719112653793,0.0176136786158341,0.00414377100664809,0.00959578409142292,0.0233729683713699
"681",0.0151341654458765,0.0184512481529386,0.00491653627317845,0.0251506955157619,0.00178428873453407,-0.000766511571019701,0.0390034272392792,0.0198071965583018,0.0102123557085469,0.0129871590421937
"682",-0.00149094854343157,-0.00076560185929897,-0.00978476150855834,-0.00536693096044405,0.0125760193290301,0.00493290766646504,-0.00488686147118778,-0.0121390267225617,-0.00570521446480976,0.000441898573175337
"683",0.000637589306714759,0.000766188454604411,0.00494062211067314,0.00282634577453944,-0.00890110376697661,-0.00534516960289633,-0.000223242202637253,0.00607192921235544,-0.00674449392971577,-0.00883775159514855
"684",-0.00253004018351544,-0.00918587027063011,-0.00983286864343946,-0.00871121762823956,0.00229823124344164,-0.000657838029681335,-0.0158518285608198,-0.0148145589403661,-0.00314175540978534,-0.0218456740229847
"685",0.005824684495918,0.0113310523457915,0.0129098771787894,0.0152495617114261,0.0020831789723359,0.00263388750417271,0.0309231485236769,0.0158730608704647,0.0133183914872064,0.0164083024803074
"686",-0.0083124692345149,-0.00789405509712859,-0.0107846517383481,-0.0150205055845773,0.00301527111446309,0.00218909426209368,-0.0335256899572114,-0.017544204065393,-0.00842777181554688,-0.022421542462665
"687",-0.0110193134215487,-0.0202770018187692,0.000991191752180764,-0.0196434787275049,0.00290200980375266,0.00273080077298093,-0.0330805035849963,-0.0181356572998509,-0.0129515225548613,-0.0128440036923365
"688",-0.00533264411545975,-0.00445378640006766,-0.00792068486179986,0.00421855260339865,0.0127137638677162,0.00402996981216597,-0.000712840745710208,-0.000852677427931936,-0.00563816487017432,-0.00789966405563647
"689",0.0179031295943288,0.0142102108393836,0.00798392299984241,0.0128643359871616,0.00877681731237967,0.00173451901191735,0.0389918232682089,0.01450478833359,0.000515494845360953,0.00889941747812428
"690",-0.00300951179012898,-0.00155657065293757,-0.020791893087561,0.002332480574605,-0.000910370662699167,-0.000431655804936981,-0.0167050168512644,-0.00616745805197239,0.00391547643744028,-0.00371406505878014
"691",-0.0038681412854874,0.0015589973424488,0.0050555198690907,0.00620677000005365,-0.000911213933313726,0.000757904547257882,-0.00698131854902306,-0.00310296657953057,0.0145745458277737,0.0279589470361863
"692",-0.0248132238370308,-0.0298389535445709,-0.0251505997569924,-0.0272425740361095,0.0136949921268299,0.00752288067971785,-0.0424187098903754,-0.0200905103144361,-0.00971167445041321,-0.00634633504819593
"693",-0.00466122473058728,-0.0090934695047592,-0.0134162634793791,0.000264159318631219,-0.00692045480046044,-0.000431289835528981,-0.00978965325916836,0.00664168744987492,0.00490350398307782,-0.0100365005487431
"694",0.01492814969728,0.0145750190693832,0.0083684591103419,0.023243884851571,0.000101317129514777,-0.000107316190027462,0.0269404601997623,0.00114770006327669,0.014740235394727,0.0322580997056205
"695",0.0143244642370375,0.0188882916403061,0.0114105614416868,0.0165203918460199,-0.00989743212641514,-0.00323449705457279,0.00024082087998889,0.0157589725096499,0.0246443498296935,-0.0120535907304756
"696",0.00274849282374334,-0.00261133209011211,0.00923101585352404,-0.00101602599426254,0.0117301739214632,0.00638198330182416,-0.00312830950708609,0.0146684089870359,0.000782186163298615,0.00180756951475836
"697",0.00765595763610905,0.0172777671948625,0.0111788800846626,0.0122014906953221,-0.0104847611780307,-0.00365428088669695,0.018827038450439,0.00917442626073139,0.0125048650595461,0.0198466927695415
"698",0.00609713271991374,-0.00643327403292349,0,0.000752991019056015,-0.0229248260457207,-0.00959997984501326,0.00971346523188754,-0.0024791726618546,-0.00771905642337956,0.00398048486315061
"699",0.00391539136864671,0.00880577961144224,0.00200982885356793,0.00828147060005624,0.00156457147691547,0.00294042543387474,-0.00164230924843101,0.00386634948692066,0.00700118658114302,0.0202642210679891
"700",-0.00204322634345577,0.0023108187218035,-0.00501507326917994,0.00174219567369316,0.0052061290521197,0.00228058406238185,-0.0150413758960652,-0.0068775481396679,0.00675940530628449,0.0112263661355538
"701",0.0172159240067151,0.0217723237007295,0.0110887303889129,0.0322977200781325,-0.0148113980227923,-0.0068260890580143,0.0367454190091967,0.034071644143266,-0.000767331656103321,0.00768576514257147
"702",0.00365946067134337,0.00777135947957297,-0.00498504333414773,-0.00553534903709207,-0.00462568832887089,-0.00327254629487972,-0.00759485856416253,-0.00482153664353502,-0.0126703685928202,0.0101693954337263
"703",-0.00747416273480284,-0.0121888881051806,-0.0180359893991748,-0.0137947722452734,0.00813255546658076,0.00459744208489288,-0.0271339976735496,-0.0156125563487228,0.00311101494156141,0.00251683053248986
"704",0.00826492779311749,0.0151095431787405,0.0163266692943511,0.019141240332518,0.00785752389880701,0.0015246631115049,0.0231230889831713,0.0210554933948945,0.0101764198488079,0.0142258758004092
"705",-0.00528313379138046,-0.00297725216753553,-0.00301226669737742,-0.0132436317111891,0.00540525673851655,0.00228445764685525,-0.0186391220958786,0.00107147373602734,-0.00777132281191617,-0.00618816184932824
"706",-0.00897330523464779,-0.00273682980731138,-0.0030210397000684,-0.0053685093597583,-0.00599612939100702,-0.00227925079494762,-0.00783481688147092,-0.0064205758857574,0.00319089157205354,0.0211707498222049
"707",0.0101641821901157,0.00998022158857981,0.00202006951088252,0.00834169645963723,-0.00488856585254904,-0.002937222411729,0.0224931175395586,0.0123856066005277,0.00163853493975918,0.00812996973268176
"708",-0.0114336987057665,-0.0170455771646074,-0.0231851606753357,-0.00827268820571991,-0.00752607555883233,-0.00490927926080964,-0.0109989275841397,-0.0250002873667224,-0.00413779838602391,-0.00362906586020384
"709",-0.0108251656885651,-0.0160845303589339,-0.00309623012421556,-0.0125119197793441,-0.0129541395659457,-0.00570069262373685,-0.00615245644881701,-0.0155479387755608,-0.0157502853560786,-0.0182111281800219
"710",-0.00458339267459684,-0.00740717810958913,-0.00414088338497987,-0.0173912557616673,0.0136572239332509,0.00860042605468903,-0.015238206513719,-0.013577464091747,-0.0000982034154898281,-0.00700753571954482
"711",-0.0188873244455258,-0.0270201215367053,-0.0103951616139117,-0.0457650400046924,0.00473691207695714,0.0030611511078904,-0.0418279768866001,-0.0410110578336438,-0.010996514698017,-0.0257368123829955
"712",0.0214537151178473,0.033060041075766,0.0157564563451238,0.0442500956981544,-0.0108950463711095,-0.00479552751742263,0.0431489935511871,0.0330987972258263,0.0194579464074871,0.0311036398292528
"713",-0.0289735006627507,-0.0358422105021725,-0.0124094065317916,-0.0466885455823985,0.0145100626277235,0.00744740925920206,-0.0191095702160147,-0.0221146264313163,-0.00155811663145167,-0.0252065640847321
"714",0.00733909242675712,0.00743482528050565,0.00942421054594011,0.0149055153049056,-0.00441948512556944,-0.0026312570967344,0.00147953295048509,0.012756816778654,0.0138495856222527,0.0173801378940006
"715",0.00316331609481613,-0.00764362494821891,-0.00103736846629121,0.00157328423189318,-0.00999520718372893,-0.00230854918018075,0.0142821076229527,-0.0031488536104165,0.0241462440831046,0.0141666878942486
"716",0.00257990762296711,0.0143422750655298,-0.00207695295902721,0.0185915585521557,-0.00913902662417798,-0.00275391843575767,-0.0179653606756314,0.0103388055061582,0.00601163823043049,-0.000821681464220014
"717",0.018394889458113,0.0172823647405238,0.00728421823616232,0.0205652587437533,0,0.000220772984202533,0.0207664322008287,0.00682188716084164,-0.00112040151485349,-0.00534540630864588
"718",0.00262045879813622,0.00205909936923998,-0.00619858270368201,-0.00125921694758158,0.000965689575745277,0.00298258920631933,-0.0154999121765528,-0.000564323557473156,0.00420636555786991,-0.0177759529768661
"719",0.0227760567203108,0.0300539828671178,0.0114345022474192,0.0368222685776973,0.00117792058898147,0.00044013576432067,0.0469864037647583,0.0364404596607244,0.00707439262775766,0.0164141340305319
"720",0.000182599183834231,-0.00274303940326082,-0.00719413924722501,-0.00462204763295937,-0.00181946942966404,0.000770585536217006,-0.00493471091817477,-0.0152630711220854,0.00184857192257004,-0.00496887633467813
"721",0.00510995021964256,0.00175038422260387,-0.00103531284679392,0.00855360277475592,0.00418137329358048,0.00285983766216447,0.0184183648257794,0.0102409557856311,0.0111633823338257,0.00665829530987594
"722",-0.010167696059034,-0.0107339744818069,-0.0165802085732625,-0.0222923300365786,-0.00181454810480819,0.000328406478833587,-0.0118246715979292,-0.0167126128432011,-0.0126824728591692,-0.0148822347476368
"723",0.00541139324468309,0.0126166249993314,0.00948357629684993,0.017100548928064,0.00459933409463686,0.00076754435171944,0.0133738413281212,0.0189468344513304,0.0141391647180407,-0.000839266802493133
"724",0.0145042732344243,0.0174436272587997,0.00939457576937519,0.0250970002103841,0.011712378039878,0.00536847101105375,0.0226903705517387,0.00929748327705671,0.0172225171719067,0.0289794580824827
"725",0.00116903630824305,-0.00612294206419506,-0.0113754093084381,-0.00356536994449264,0.0053670038750675,0.00217953476714094,-0.0142627426510116,-0.00623132005983107,0.00304581213954513,0.00489801833895021
"726",-0.000628859559538952,0.000739276935530553,-0.0104600316042904,-0.00787185040250526,-0.0058620006386072,-0.00250109941940069,0.0165363812565711,-0.0073608536560843,0.00250066086897682,0.000812252937989699
"727",-0.013031443104266,-0.017729907423624,-0.0232560724859066,-0.0185142917507549,0.00179004300345365,0.00119909681008412,-0.0198824735619541,-0.0192258971422326,0.000445461024498828,-0.0142044773407461
"728",-0.00355124053682887,-0.0127847958992523,0.0075759356103664,-0.00416467141582033,-0.000210198656862892,-0.000109453824059469,-0.00760766069543639,-0.00588057837740419,0.00569901142389106,-0.00123505925958234
"729",0.0127024224739125,0.0210763573545223,0.0107409754289889,0.0209102893704922,-0.0012617405967531,-0.00141518795656548,0.0113826873151355,0.00957716279652421,0.0119532404470826,0.00453423541191289
"730",0.00153387267892646,0,-0.0127522813059359,-0.0055419869794564,0.00631626139365316,0.0051252824055712,-0.0146995740985699,-0.00809113763026559,0.00384987309607254,-0.0114896742436308
"731",0.00351398282673587,0.012683456597038,0.0172227125925397,0.0116306421360035,0.00460207555651237,0.00336271237435271,0.00396287491369396,0.00759492856908883,0.0164734589957258,0.0240763949254048
"732",-0.0162507676880993,-0.0348723632082344,-0.00846549375390604,-0.0388022500777868,0.00374875179541623,0.00454100474460817,-0.028325938422083,-0.0304299818393655,-0.0133768218133213,-0.0113497883869876
"733",0.00337710415460601,0.000763562798468342,0.0202773860030345,0.00971815601307213,0.00238615044996027,0.00161500397374326,0.0375151354995864,0.0129571531205996,0.00504085703182455,0.0110701708064096
"734",0.0123700657685928,0.0218658584955829,0.0345189874417955,0.0286279116012986,-0.0111395868200357,-0.00551562301008801,0.012897016552837,0.0264353902117527,0.0150466794798225,0.00729925362220607
"735",-0.000448914070415918,0.00273737068944824,-0.00404425414547505,0.0040786204486214,0.000839610314814943,-0.00205692704926219,0.0147794906372876,0.00138474089523455,0.0153348359686873,-0.00684387248095841
"736",-0.00782065945029065,-0.00719610875508869,0.0142128641795316,-0.00931907692848499,-0.0103853067077385,-0.00466561548632327,-0.00851466124722944,-0.00940265402041207,-0.00402754656821624,-0.000810606791958768
"737",0.00570780874868726,-0.000249891099231458,0,0.0091655206369412,-0.0105998472777674,-0.00741423958641096,0.026892741991245,-0.00111674140859985,-0.0417017449461267,-0.00811360440726594
"738",-0.00153159229843058,-0.0059999383862267,-0.00800778021670656,-0.00860434041937763,0.00128600808231094,0.00274545333741427,-0.0173856931743613,-0.00475148209284437,-0.00562636483516488,-0.00899800029003262
"739",-0.0110966778077376,-0.022384451885612,0.00302701640766601,-0.018562946841339,0.0014975241733246,0.00350599953803266,-0.00604700220548415,-0.0235885209362284,-0.0190964899735082,-0.00990506872576724
"740",0.00374040611327664,-0.00128648472749404,0.00301811965563337,0.00614088718748018,-0.0045941101829704,-0.00196526096249516,-0.00135168208266068,0.0115040865448945,-0.000991446624374337,-0.0125052544077175
"741",0.00563534411920186,0.00154593827397309,-0.00802399243475138,0.00585966856992859,-0.0114843316745906,-0.00339029275377511,-0.00293339599609366,-0.0062555934671148,-0.000180404192724803,-0.00548755975720583
"742",0.00424796226575941,0.00360039837704096,0.00606687545370455,0.00364044536519725,-0.000108325643666918,-0.00493843946340544,0.0144831926594713,-0.00457775283864992,-0.0135354629128316,0.00509348414873867
"743",0.00684013906992131,0.0112762317626263,0.00100501863241287,0.00677175256601892,0.00119455716391959,0,0.0194065718869671,0.0091981234140337,0.00841564215148205,0.00548978970308478
"744",-0.00464839078762613,-0.0114036637998782,-0.00803225513145811,-0.0103290474067261,-0.00444699944339066,-0.00319869779055482,-0.00919065521711471,-0.00882922908521222,-0.000272124460669931,-0.00461984469599885
"745",0.00152699338544315,0.0110227180631797,0.0151820901828867,0.00582511066802516,-0.00119802218131815,0,0.00596296584584133,0.003735197863308,0.0125215226614783,0.01729955854448
"746",-0.0120160770071296,-0.0268762398686789,-0.013958038636013,-0.0287161412075658,0.0164704487057412,0.00885222045735978,-0.00636618329345118,-0.016031921908676,-0.0380858513517646,-0.0153464185073455
"747",0.00565744106568777,0.000260716399815619,-0.0020223517252338,0.00273258219633177,-0.00429279787660941,-0.00493570615755068,0.00773283100543543,-0.00212822530161971,0.0149990782559746,0.00421237281712639
"748",0.0101622662276957,0.00763783109209304,-0.00303928469283254,-0.00123837892240031,-0.0177819966304478,-0.0102502916435853,0.0120585371572226,0.00207345286714311,-0.0183570450213046,-0.00964764890606939
"749",0.00359334441044479,0.00833551411023814,0.00799825554569611,0.0100778107474988,-0.00559548080200289,-0.00445448877524535,0.010615591839146,-0.00443395688130888,-0.00729311848414538,0.00720032777982405
"750",0.00196885524023593,0.0105915094602502,0.00305180825313744,0.0099032295628938,0.000220180031544004,-0.000447457323446199,0.011289275621158,0.0142518019299194,0.00357921265101657,0.0176619629297825
"751",0.00473439321118052,0.00255648387632901,0.00709951822549604,0.0100518715819369,-0.0103695799441418,-0.00358087089704118,0.0126419915583631,0.0014638277479655,0.0169873106432479,0.00578508727199134
"752",0.00213355642018986,0.00484425611228545,-0.00402827723722377,0.00339806273985888,-0.00278673191099676,-0.00269510893392111,0.00359719499374811,0.0055535308575283,0.00175343298492603,0.017666362905564
"753",-0.0014193644975462,-0.00126837402613045,0.00404456988603008,-0.00358103759363482,0.00659634602661119,0.00263947606231918,-0.0143369274446585,0.00784913471453708,-0.00994935025473931,-0.00201862644316708
"754",-0.000355241799199435,-0.00152468063938893,-0.0110777476192624,0.00437122252819178,0.00657576127771931,0.001800520754901,0.00171167484375734,0.00490331494514185,-0.00502466730227336,-0.00121349249101033
"755",-0.0095984419753169,-0.00865119742805986,-0.00814677280124576,0.0033848575967228,-0.00476178409074846,-0.00482978996155325,-0.0194325369886398,0.00143510573087591,0.00355370803329258,-0.0028351171688914
"756",0.0169599699359422,0.0266936992362803,0.0256674617980064,0.0291567302181714,-0.000889805891861051,0.00248300584642402,-0.00239518953968643,0.0214965938818512,0.0232038490952167,0.0251827673620635
"757",0.00264679089558406,0.00100022463171712,0.00600600891839354,0.00725800446594493,0.0064579601878394,0.00439166183284567,0.0024009402466505,0.0103811326571508,-0.000910801432309705,0.00118857325538912
"758",0.000704117811222371,0.0012487199879283,0.00398006247005456,0.00209191616582083,-0.0133861585788294,-0.00403605213348246,-0.000435445375123078,-0.00527612771652297,0.0164995902415568,0.0178076370356166
"759",0.00422160461686216,-0.00324258248158593,-0.00891945070094546,-0.00579895417318466,0.00168218444208179,0,0.00893223152136158,-0.00670000440234397,-0.00618780367343197,-0.0124417099344923
"760",0.00332760743166505,0.00800774607708243,0.011999768061989,0.0079326185826214,-0.000447924137659816,0.00123807254140762,-0.00669378556484057,0.00533969254300337,0.00496303013896404,-0.000787390854466552
"761",0.00139653116730631,0.00819274230483069,0.00889332836314916,-0.00208331425862884,-0.00548730597867286,0.000674705856663183,0.00478259050304541,0.00419347991402996,0.0132889912914882,-0.00315212641401641
"762",-0.00932662174766974,-0.0137894159758014,0.00685614624482267,-0.0160056966003524,0.0171172427304269,0.00718924562637402,-0.0168758601556951,-0.0105787928459463,-0.0209127163653118,-0.0213438275954736
"763",0.00844676316529891,0.0114855414687436,0.00583626349818367,0.00306481943066061,-0.0116259471029098,-0.00479563034048969,0.0187063319710978,0.008160024629706,0.00950314977831757,0.000807826564948932
"764",0.00270416567113529,0.00049353307909783,0.0145069065228649,-0.00258528254177159,0.0140032409882518,0.00470641963337681,-0.00345673300514737,-0.000279375069273335,0.00439302488440885,-0.0052461774260445
"765",-0.0112240892936356,-0.0180115917073583,-0.00190639202344189,-0.0115455410711589,0.0061862906010044,0.00446204766177427,-0.00910437983349965,-0.0117252040182162,-0.0104436134110829,-0.0113589960663488
"766",0.0124958550612879,0.010553085537429,-0.000955226957606747,0.0202619621270319,-0.00285508662072376,-0.00177680216380705,0.0199077169259276,0.0155366332412985,0.00595341867261934,0.00656544367339817
"767",-0.0101689194968066,-0.0256091049171847,-0.0219885040304547,-0.0240653390219069,0.0101296530948318,0.00344833788952315,-0.0102961980560727,-0.0255910462561425,-0.0231348194889208,-0.0187525843160991
"768",-0.0192289934796976,-0.0308752948201553,0.00488766874068824,-0.0301651491827765,0.00457825828551561,0.00365913844763766,-0.0283915892048558,-0.0191264898650184,-0.0144115932731488,-0.0124636054323451
"769",-0.0222919842308903,-0.0234332398756725,-0.0107005589623003,-0.0222167748865835,-0.00173609726039203,0.000882962834260814,-0.0229757186628876,-0.0189173025533824,-0.00186276422102727,-0.010517487817516
"770",0.00512809280584769,0.017524716338303,0.00786651767064472,0.00732146828419844,-0.00456533375692769,-0.00220713314730414,0.00730592360452276,0.0201719109365717,0.00289264725002591,0.00467680669095438
"771",-0.00419074326284985,-0.00370958512896236,-0.0107315618377523,-0.0208021174646518,0.000328468266091786,0.00199092654701882,-0.008612632515968,-0.013666798213687,0.000744277984435771,-0.0110028558895792
"772",0.004757338147928,0.00505333073230063,-0.00591750772388244,-0.00255930991795517,-0.000545966247105234,-0.00231793804831659,0.00914503886797724,-0.00353775375647924,-0.00957604145734536,-0.0145486749141351
"773",-0.0114722728321875,-0.0254037503961766,-0.00992057129367541,-0.00692831000319472,-0.000546264489078241,-0.000332478928401936,-0.00951540308745791,-0.00562110494651935,-0.000469313812722416,-0.00347368256874803
"774",-0.0108688192321506,-0.0119467194937515,-0.0140279828912674,-0.0108530775311385,0.00874152575537535,0.00387472691152313,-0.00663323917673864,-0.00684319996526905,-0.00488358363400876,-0.0113289556147773
"775",0.0155508149936547,0.0200604299099711,0.0101623261829851,0.0269071034388702,-0.00907698218593589,-0.00342957260840804,0.0181903116991693,0.0161771673291002,0.0225556721645497,0.0242397840215776
"776",0.0121030626146383,0.0161638260999319,0.0191149402585016,0.00814069925838501,0.00285267474256146,0.00166524091296005,0.0165084797844555,0.0232901431266539,0.00719888338161301,0.0215144674378465
"777",-0.00498219051431548,-0.00954418493789488,-0.00987186472326829,-0.0058038537165821,-0.0115962409099601,-0.00476580756582645,-0.0115682769145561,-0.0149811290518801,-0.00394025485036897,-0.0122155473463933
"778",-0.0308663043719247,-0.0455032754197587,-0.0189429510840941,-0.045177717775055,0.0158269716854453,0.00824010071730741,-0.0373627669530265,-0.026616184834914,-0.0398343525253271,-0.0332622435452573
"779",0.00206704154292514,-0.0190687707164856,-0.00203268006032953,-0.0111640947781537,0.00217902460276487,0.00320230269757182,0.0187049997888982,0.0012020172337206,0.00297017333610694,-0.0127923788437495
"780",-0.00721926119537286,-0.0111490041287868,-0.00712807864379894,-0.00994619072955283,0.00130465621967657,-0.000880053448209406,-0.0227217176863455,-0.0237092153020096,-0.00611386129155522,0.000446913439102747
"781",0.0125602848668471,0.0361372096244117,0.00615372709546302,0.0325817030878084,-0.00998852508750958,-0.00539920909268121,-0.00305349843826097,0.0230552633824541,0.0131680410114567,0.0178651962283896
"782",-0.00195874459579204,-0.00530114778069601,0,-0.00262929923229971,-0.0095421363477225,-0.00276938275985306,0.000706854334150187,-0.00120170028784505,-0.00275117151119741,0.00394900110499585
"783",0.0104666848928514,0.00729300609233108,0.00509680679755409,0.0263641908979255,-0.00542517370029616,-0.00122180612530676,0.00870972916738588,0.0072200930741857,0.0191209469428955,0.0118007183910438
"784",-0.000832509046514218,-0.00863261356588541,-0.00608528432121891,-0.0125866675613472,0.00411884092398473,0.00233562407503296,0.00910175074287745,-0.00627243272250777,-0.000840063497808186,-0.00561547411050289
"785",0.0157344334022673,0.0230339367713766,0.0102043760199531,0.0257545402558237,0.0018845209681404,0.0022192291249159,0.0268268847187101,0.013526189445807,0.0241031574728778,0.0304082808699191
"786",0.00473921445974002,-0.0010984699388491,0,0.00355091390665807,-0.0113983839360217,-0.00531460025148778,0.00945975237064656,0.00207559856322193,-0.00337532375364014,-0.00505895277612167
"787",0.00589500285245648,0.00494793902956681,0.00201988605115533,0.00379039259428104,-0.00403007671831268,-0.00356191929361616,0.0133865890210627,0.00562276722828958,0.00668194965675051,0.0088981828450192
"788",0.00207366809391529,-0.000547150216263725,-0.0161288823685576,-0.008559782149268,0.00539450361079319,0.000558785409576545,-0.00021990918960324,-0.00971154065534863,-0.00463722482349815,0.00588001847142516
"789",0.000180061645440155,0.00136843988333069,0.0122948455093081,0.00126958127691945,-0.00413543489606805,-0.000781422893601169,0.00418388529695335,0.00267470923632263,-0.00365397822550495,-0.00542802922543661
"790",-0.012144750352543,-0.021044364453649,-0.00404830797403222,-0.0230788310137293,0.0156036500832322,0.00759736827008117,-0.00789459888361199,-0.00859504230411057,-0.0108187494269734,-0.0163728741687471
"791",0.009197602825606,0.00949236176100743,0.00203244136729341,0.00960535689209152,0.0024310484313268,0.000555217835431998,0.00972616078761002,0.00956642279359055,-0.00491239229689866,0.00810937083926322
"792",-0.00135354717961234,-0.00884997593814207,0.00202819982355273,-0.00822852086455317,0.00562473630806548,0.00365640488641827,0.00503420277481359,-0.00444183391804687,0.00884870520819003,-0.0169348735900949
"793",0.000632342747397763,0.00502267857430394,0.0060728779828314,0.0101115964513554,0.00515316876923677,0.00154607608764201,-0.00239561616387718,0.00832808558716258,0.010340707420196,0.0176571726432413
"794",0.0103850706189417,0.00222073788719723,0.0100605352912233,0.0169405601670971,-0.000437835962671329,0.00103938759169475,0.0102620714310853,0.00855489321098246,0,-0.010156572821003
"795",0.00277024348478849,0.0132963968227231,0.0029880051395057,0.0113579192271078,-0.00131374825710096,0.000552198224127665,0.000432564326557916,0.0152089766944872,0.0145298090103263,0.0106884025606933
"796",0.000891288189557748,0.0120285887147396,0.00695169841061216,0.00124778082010479,-0.00252137120592644,-0.000993310067738729,-0.002160648574831,-0.00316914830177673,0.00549450564297893,0.00972926960187404
"797",0.00302762441988014,0.00135080601102855,-0.00986224263689717,-0.00523432036513605,0.00527489957080252,0.00176708075810073,0.00411345663736173,-0.00115605826253162,-0.00716648769595518,-0.00879774891871954
"798",0.0142934478037138,0.0207712515141878,0.00996047526069699,0.0260584601525413,-0.0131189760499506,-0.00474156786714153,0.0228547460751847,0.0205440001595214,-0.000180492643138241,0.0118343758967849
"799",0.000175235467013257,-0.00396424532497763,0.00690301103588853,0.000732784668097564,-0.00520610664118448,-0.00266017352124348,0.0124367980483882,-0.00482015063712171,-0.00839275351308999,-0.00125311570013642
"800",0.00166235949577187,-0.00159163003865337,-0.0039177773146245,0.00561232844428261,0.000222421609271217,0.00255604177528457,0.00333119959619599,-0.00113908952773878,-0.00145609760073084,-0.0108741776279682
"801",0.00445582024654612,0.00425194903093185,-0.00688291066840896,0.00703750822108073,-0.0025606566172347,-0.00166308556584605,0.00539569173369903,-0.00912767121710589,-0.011392635696385,0.00295987758725458
"802",0.00417501786181473,0.00846767893522582,0.00990095527429835,0.0002405887860506,0.00368392047826749,-0.000887916197431782,0.00495351218788964,0.00690880215177558,0.00119846039274951,-0.00252956316850506
"803",0.0000867070301300288,0.00472336337267065,0.00980397377413267,-0.00337250883304729,0.00622709708485925,0.00155601325128063,0.00739310059961085,0.000571573771312339,-0.00598527635332002,-0.00591707919774553
"804",0.000259864445077751,-0.0107077904377365,-0.00485422350566778,-0.00725166379920117,-0.00132701484793685,0,-0.00285435926033017,0.00171459566638665,0.00379809181467605,-0.0119047301272583
"805",0.00796618754936551,0.0163672507196191,0.0097559470795805,0.0129047543699248,0.00796879692332975,0.00388265331861914,0.0259665664865298,0.0168279889644607,0.0188261441599655,0.0133390202979642
"806",0.00592722910305654,0.00285744304183155,0.00386489652255761,0.0108176527007284,0.00428192281470441,0.00121564435704036,0.0121558032270168,-0.00112230467995478,-0.00733701073664839,0.00891716287918798
"807",-0.000512366055897773,-0.00699318721859388,-0.00673736658287649,-0.00761001008139306,-0.00327900591364783,-0.00264899047634015,-0.00393744864043344,-0.00224639080634093,0.00684369036750399,-0.00210443502469138
"808",-0.00506187785209156,-0.0112152590656338,-0.00193802308956659,-0.012940768814997,0.000986454965333561,-0.00132773969291022,-0.00849967009816088,-0.0161985735664228,-0.0186695402816581,-0.01223100333295
"809",0.00534600883040892,0.001318880022535,0.00485436602627876,0.0036418868864192,0.00109603696659755,0.00332435099976047,0.0103666215781821,0.00660926030732645,-0.00489470820922344,0
"810",0.00703345306182768,0.0057955067675397,0.00966177326044404,0.00701507820353475,-0.0047070505824357,-0.00209878653772022,-0.002761975562251,-0.00256972718282922,0.00529002320185601,-0.00426988417232754
"811",-0.00485476629399162,-0.015453061419083,-0.0162678046629511,-0.0148931309743677,-0.018255815826493,-0.00996176251052405,0.00316567218357044,-0.0151685526087474,-0.0186484213441653,-0.0111492962624892
"812",-0.00162647812561278,0.000531870858254679,-0.00583677757054313,-0.00268227428688317,-0.00638432984960113,-0.00368890841896541,0.00157356658525654,-0.000871806233994521,0.00451548435045668,-0.0056373907344931
"813",-0.000599689393745106,0.00771089579266704,0.0156557480326001,0.00489004707387708,0.00281761349639664,0.00235665778002381,-0.0035799701874587,0.0116347180234253,0.0169507119025165,0.0017444157174622
"814",0.00634751423248803,0.00949846350947969,0.0125238674678441,0.0180047235147143,-0.00382213353333105,-0.00145511027601164,0.00439095891827868,0.0212762499097334,0.00147346906615597,0.0226382280421098
"815",0.000681719206399922,-0.00444314396469414,0.00570907535511278,0.00382405962527943,0.00315962615834664,0.00100826288050282,-0.0019869835031161,-0.00281489628905429,-0.00717240459770119,0.0021286238789695
"816",-0.00340709723494648,0.00656334430982186,-0.0122989679906186,0.00285706758457405,0.00686320593197642,0.00235247590243826,-0.00895870615528405,-0.009599156097294,0.00907655821916675,-0.000849649729898538
"817",0.00683765778424972,0.0164320700112832,0.0153256100522006,0.0261160851349849,-0.00244485018369733,-0.00207335869283443,0.00462021004127644,0.0193839868020693,0.0120239103815671,0.0195577740490089
"818",0.00814952009045267,0.00538857674873583,-0.00283012055931375,0.00902338252970147,-0.0166390011557024,-0.0089825008745642,0.020795450071841,0.00531351885392772,0.00571374014667625,0.0158465370998924
"819",0.00235758047230705,-0.00689110605000043,0.00283815287411326,0.00298104710006952,0.00160146656698767,0.00294605687855665,0.0201767568028097,-0.000556663895843079,0.00126251241106057,-0.000821006858102935
"820",-0.00571235751315702,-0.0110513790365541,0,-0.00868772932427742,0.01278339621244,0.00621296073131439,-0.0215056392221097,-0.0158638201144654,0.0131495903192793,-0.00369756658899045
"821",0.00346393887988072,-0.00051949932262918,0.00094342891457555,0.0034594250940474,0.000450494394407697,-0.00112207962426714,0.000392249815246881,0.00735282362038792,0.00142238423721897,-0.00164954680753537
"822",0.00656732639124091,0.0145605882389443,0.00282745305834364,0.00620561099357175,0.00236594543575563,0.00112334010130599,0.0158890937709739,0.0106680173172986,0.00878825550309359,0.00206531912904606
"823",0.00158944498164293,0.00794463764430087,-0.00187973685174114,-0.00799437436875938,0.00528175504573447,0.00269504630564876,-0.0065649742858237,-0.000555356089336212,-0.0055437962473055,-0.000824475860280893
"824",0.000751679231047575,0.000508306057635632,-0.00188316633578989,-0.00207270612176458,0.0032424817892851,0.00190295035927446,0.0227403854312205,0.000555664681100465,-0.00283160777220404,0.00371290560147886
"825",0.0113492407261597,0.0142310267852936,0.00471717227028035,0.0147670930014832,-0.00702064036395078,-0.00268227073315264,0.000950144973224543,0.0127778573211788,0.00301709995532695,0.011508480076293
"826",0.000825169331444497,-0.00350765076656656,0.00469472178742358,-0.00545702221329536,0.00112182773438585,0.00168160431393161,-0.0248719140725484,0.000548541375342548,0.00548529598766079,0.00365708345691451
"827",-0.0159122450692011,-0.0213729377627793,-0.0186915215990745,-0.029263670887702,0.00728712630516259,0.00604061658716204,-0.0208329059942872,-0.021655769262416,-0.0212054901679632,-0.0182186646443475
"828",0.0037702695579851,-0.00385417157812096,-0.00190510723868609,-0.00400389181650895,-0.00244841192388989,-0.00244592357326467,0.00377753607045817,-0.00504338414739547,-0.000809025544930342,-0.0127835421184697
"829",0.00893052706465536,0.008511865875104,-0.0038165347050455,0.0118233141379931,0.00356951229568248,0.000445253259024003,0.0156499734788473,0.00816691082409826,0.0027889968009176,0.00793648541716063
"830",-0.00181992092845296,-0.00818408429080242,0.00383115644658427,-0.00327173910195155,0.00822587687098708,0.0032315049101963,0.01872436449549,0.00139621958355507,0.00762604528643496,0.0049731226595251
"831",0.00298370060646258,-0.0108302006462316,-0.00858741319550471,0.00422027173815365,-0.00297716914754609,-0.00233229317252581,0.0145509691930612,-0.00223130527550597,-0.00418486339924962,0.00247419288560891
"832",0.00652776468099248,0.00860234775197388,0.00673705575356642,0.00537008119075999,-0.00353843377902752,-0.00278303490489817,0.0130214040656007,0.00698930302885303,0.0120708695304317,0.00658156363703033
"833",-0.00377626986444479,-0.00155042239243597,0.00669216804480621,0,0.00110993715577656,0.000669695070709242,0.00633385874685577,-0.00111053250799054,-0.0038872867941111,-0.00490381329421719
"834",-0.0236507170806401,-0.0445251968288469,-0.0180438918226914,-0.0357642987186685,0.0140780991519707,0.0093711191558894,-0.0316548883812684,-0.033074039363611,0.0166740310421287,-0.0151951590075315
"835",0.00759606076559471,-0.00487681780195393,-0.00386823771795131,0.00842976018437747,-0.00852636868848033,-0.00508440058960269,0.00344108738394722,0.00632385034154548,-0.00279158168345772,0.00333606789495611
"836",0.0123972045889835,0.0185136715417491,0.0116504898647181,0.0164793293259931,0.00419002334158702,0.0016667046867922,0.041341033231008,0.0159953815271785,-0.000262435487051516,0.00789703081839277
"837",-0.0169615826357477,-0.0155039502880563,-0.00287892480919649,-0.0119825599885814,0.011527989540324,0.00609937865321708,-0.0311012555203097,-0.00590382169419268,0.00945049010719701,0.00783502902155764
"838",0.0129619496815805,0.00705974798501985,0.00288723694727411,0.00546936966620049,-0.00130720390974026,-0.00262074422368219,0.0309665687315039,0.015271549849001,0.00320736821075451,0.00490995854541798
"839",-0.0235147970547508,-0.040172792615417,-0.030710193673815,-0.0458844541926453,0.017995124232111,0.00676201567029056,-0.0234429150767783,-0.0406688275193382,-0.0074310894124836,-0.0268729322961048
"840",-0.0059562981654534,-0.0269661730644521,-0.000990220522241292,-0.018096332395873,0.00589244981508941,0.0038537331566777,-0.0140661029305693,-0.0153889694463277,0.0019151475080923,-0.0225941773588147
"841",-0.0332136953596536,-0.0534063745849577,-0.00594648475066284,-0.0408985736986154,0.0308878545842948,0.0109690223374803,-0.0401370247383079,-0.055145962599076,0.0295421158933744,-0.0196918202787819
"842",-0.0148751011527959,-0.00579460813889987,-0.00897312934889394,0.00526410105838915,-0.0125015032635404,-0.00271275859605202,-0.0168452164621952,0.00530584657532529,-0.00185670523852988,-0.00524014825566066
"843",0.0440411111528629,0.0763806686291064,0.0281690793975469,0.0720088067259339,-0.0207162363023378,-0.00761523106606388,0.0659140513623619,0.0509156729119604,-0.0059186354760794,0.0193151962987981
"844",-0.00284084828624931,-0.00541487246494265,-0.0225048702743458,-0.0180751801445852,-0.00256387548630566,0.00120574168064946,0.0011346288147398,-0.0141802871403185,0.0262822488730119,-0.00172262936785217
"845",0.0139859231285904,0.0163323634119208,0.00900905746054681,0.0124377927983708,-0.00760454353399553,-0.00251825815833462,0.016245231950347,0.0107884048551468,0.00613291874248567,0.00819678682120339
"846",-0.0124306689352295,-0.0219903888103642,-0.00793631722899968,-0.00933679085234274,0.00658400652349145,0.00274420387167695,-0.013197221675123,-0.0103765546476146,-0.00691930795849582,-0.00855803888595574
"847",-0.0181052493004612,-0.0302683023752672,-0.00700000660582956,-0.0205852469488547,0.0173703942607437,0.00645924653878849,-0.0308907446609887,-0.0170759647891269,-0.00157593731877792,-0.0254639689982534
"848",0.000526773849757411,-0.000594243009317763,-0.00201425688343382,-0.00607770205187574,-0.0036886198776821,-0.00217612444049986,-0.00155490443409934,-0.000304915682492024,-0.00839081145491039,-0.0283436440301731
"849",-0.0136021081850354,-0.0190366680980132,-0.0171545693534733,-0.020891418944602,0.0153389274157647,0.00730405391954547,-0.0255013041167076,-0.0216464919465648,0.00108911694797986,-0.00136734681240436
"850",-0.0056940327600834,0.0042452354245881,0.00718710874425832,-0.00962813961562337,0.00333380441957787,0.000865528232914414,-0.00839027823341265,-0.00218104548267128,-0.0239350660964945,-0.00912836160459607
"851",-0.0377596094533408,-0.0314009313732075,-0.0152903306090388,-0.0496584022719958,0.021080165001824,0.0097304718017257,-0.0483478482836925,-0.0371644482944768,-0.006773566152111,-0.0207277302351985
"852",0.0145993222788321,0.019950189148588,0.00931669562067139,0.0323471575632721,0.00101709680616202,0.000535390606578368,0.0323875813798629,0.0204345984758341,-0.00535216696658036,0.010348075457902
"853",-0.0128313223687621,-0.0259782093997425,-0.0133333413632113,-0.0104443148455609,-0.00345403309904824,0,-0.0200942999739051,-0.017164387563434,0.0140600155002604,-0.000931085981564328
"854",0.00102136026880939,-0.0015687922664519,-0.00623725184803015,-0.0108253649208395,0.00489302799525171,0.0034248713938223,0.0104625278537371,-0.00840888864938694,0.00445057358612022,-0.00792165449983961
"855",-0.00602845949252495,-0.014142120283278,-0.0125523994260697,-0.000547456439640603,-0.00284024326719023,-0.00202644481601377,-0.00393444170109847,-0.00913239324315129,0.00945807762902118,0.0108030940099144
"856",0.0334982127785108,0.0621614750390327,0.0243645090436448,0.0604983506426329,-0.0226881008264839,-0.00951171249939575,0.0542616576658688,0.0513493868136194,0.00185701863883669,0.0292750765132741
"857",-0.0125497345104861,-0.0204083325621176,-0.0165457431973528,-0.0165201900906149,0.0045806167777267,0.00453174121136879,-0.0149868695841536,-0.0159672123817284,0.00160076667620235,-0.00857780778638462
"858",-0.0168237153886485,-0.0119483317127077,-0.0031547445613318,-0.0183728243722889,0.00702867989203737,0.00129279976005403,-0.0194194603553276,-0.0104998430478028,0.00866425829401729,-0.0186703822178462
"859",0.0260394633972001,0.0310078951893658,0.00527410355352798,0.0350268138059711,-0.0094997040278807,-0.00570180942599507,0.0220498915236971,0.0369776394405943,-0.00108418810493904,0.012065039772875
"860",0.00344419750082903,-0.00210542100897915,-0.00209830838654534,-0.00361699156511697,-0.00729666815707264,-0.00140620804978286,-0.00259692928612232,-0.00279091652350549,-0.015194523419557,0.00550208235748162
"861",-0.035137034100338,-0.0491259611469024,-0.0189275412089821,-0.0355194771858049,0.0268822483629039,0.0138680502459616,-0.0542757974894392,-0.0407336055579226,0.0104272889998924,-0.0310077024594181
"862",-0.0124508163597452,-0.00919188790378944,-0.0160775371012098,-0.0155914755113348,0.00766972445104286,0.00406044252371296,-0.00508276581842149,-0.00842802701507328,0.0192968869989614,0.00188232704909397
"863",0.0107119985764488,0.0111964401340843,0.00980397612574513,0.0229381830251052,-0.00497234380053801,-0.00308663482597304,0.0174541539748501,0.011768789729435,-0.00403323736987793,0.00798490818368358
"864",-0.00534589925079199,-0.00284697569615877,0.001079197993892,-0.00533894241902411,-0.00112196837929457,0.000106927991110783,0.00502084983603512,0.00387718569543427,-0.00363638016528933,0.0046598644724829
"865",0.0292314370768085,0.0491750017891455,0.0172409603913486,0.0348899934726337,-0.0178676448471382,-0.00928688890921103,0.0418402288144331,0.037978691648781,-0.0131884292167954,0.0166975025710112
"866",0.00485569051755297,0.00332625953101062,-0.00211856236203622,0.00518654209489866,0.0126825188812942,0.0063571925833743,0.0103895027046856,0.00186023112192668,0.00874170792013351,0.00136868840960847
"867",-0.00155000855562959,0.00693182699723516,0.00636955459556554,0.000258009697426065,-0.00513313156294837,-0.00085676878813512,0.0118644608659049,0.00185715627576788,-0.00341641524178959,0.00273344776777806
"868",0.0227375302925741,0.0359174215421394,0.017932552893561,0.0301778224958333,-0.00412714992512409,-0.00310740999383041,0.0216927402902385,0.0299658292513678,0.0116220737729444,0.0168104514110876
"869",-0.000357214337308953,-0.00953472624082718,0.00414503843687863,0,0.00569900377127541,0.00279498742733542,-0.00726847039784262,-0.00419880815646967,-0.00545496331027306,0.00223419928982249
"870",0.00160781490386763,0.00554250645363163,-0.00206411550078445,-0.00500758596132256,0.00813890240826365,0.0047163924007283,0.00154131058053064,0.00030117569756194,0.0130474526211677,0.000445917171275401
"871",0.00108422713179857,0.00116029864302614,0.0020683848860894,0.00452961779429417,-0.00163495768106248,-0.00202722066144789,-0.00288564284279202,-0.00671319984018726,0.00762920414062007,-0.00178259847966811
"872",-0.00286407989094339,-0.00663017906918228,0.00722394977526997,0.0172847094756481,-0.00286633311115247,-0.000748305223267853,-0.00713889817389846,0.00214078113786553,-0.0198648779636101,-0.00401780231396276
"873",-0.0165156716603805,-0.00923719139352008,-0.0122951764024348,-0.0192072068890259,0.0119084976664696,0.00599110826920479,-0.0281770259814726,-0.00762878478313433,0.00880470146029322,-0.00224111676075323
"874",-0.00310326177231335,0.0066164535159694,-0.00428386140741832,0.00257788552937188,0.00679743019423751,0.00372191171304648,0.000599711518130208,0.00491987018064433,-0.0041169206451277,-0.0166218384377776
"875",-0.0165703106565214,-0.0179265481577885,-0.00314776700412955,-0.0176454599024565,-0.00594529630244345,-0.000847081291268093,-0.0205998743428165,-0.0140756962804871,0.00289380743018963,0.00228421090344666
"876",0.00418931182652216,0.00212961180805338,0.00421054156052691,0.0118038583389997,0.00405446001676824,0.00159007366167629,0.0255194438474107,0.0117937028991895,0.0120362651598616,0.0182315253844831
"877",-0.00315208876553608,-0.00394642836892301,-0.011530485726978,-0.00684730036512371,0.00938948162768161,0.0070934586895941,-0.0114385964384034,-0.00797549081437754,-0.0136038283870344,-0.0107431451285394
"878",-0.0308751417424791,-0.0374887067849086,-0.0243903185412713,-0.0406030022892193,0.0109017647555332,0.00431071711488862,-0.0320745926453134,-0.028138342226564,0.00148650595380317,-0.0276017606022768
"879",-0.00950004931217696,-0.0072830840782897,0,-0.00665414148962507,0.00672815967207763,0.00146543475139072,-0.00985738631348798,-0.0082722161589136,0.00338091044893818,0.00372261089084946
"880",-0.00445661928332719,0.0169060250784767,0.00326092938562783,0.00723459720311048,0.00157702588096331,-0.000440098309702708,-0.0019065299468124,0.0134740030675486,-0.0381327991452992,-0.0152989615223466
"881",-0.00544937939710488,-0.00470516649971142,0.00433352107082263,0.00425655284380433,-0.00797246778214111,-0.00178189066553003,-0.0190999722884413,-0.00158203584973959,0.0123889011244966,-0.00188311652441298
"882",0.00655583288242356,0.0226916083984157,0.0204968228100859,0.0185429888066762,0.00823531925442267,0.00241545971197121,-0.0194718847475225,0.0117305664686349,-0.0167102374328676,0.00283005256186408
"883",0.0314958140304602,0.0354390152915267,0.0190272695602574,0.0221064645724192,-0.0117102369539831,-0.00314329663510859,0.0476607172103847,0.0363521758434675,0.0104712125916879,0.0225775443640059
"884",0.00989573812940625,0.0104166372031849,0.0020746355984862,0.00483491825883386,-0.00637236489753645,-0.00241791792275692,0.0107413330114958,0.000302718967200466,-0.00441691995879756,0.00919974372801868
"885",0.00746519861487882,0.00147276103581295,-0.00621114188999805,0.0121550159360397,-0.00571210088865581,-0.00263353392096033,0.0131273852938809,0.000302312665668047,0.00981146668212163,0.00182312908320581
"886",0.000648433512182578,-0.00264699371596189,-0.00520854904171719,-0.00800604073706124,-0.000403242989956198,0.00168980478253578,0.00370262966733237,0.000906559035895427,-0.00861781844695997,-0.0113739613018505
"887",0.0150886397859122,0.0253612520560453,0.00523582006731149,0.011601236223721,-0.00857058401596389,-0.00495626523932413,0.0219262326462457,0.0132849071739107,0.00869273082300093,0.0161067811886209
"888",-0.0000914130346391095,0.0025882985444825,0.00729137353099185,-0.00199433399059357,0.0100681453638751,0.00498095215937044,-0.00581500467981011,0.00327756675693869,-0.000506911114338315,-0.00181156937638549
"889",0.000273753317121095,0.0100401331944506,-0.00827279970292638,-0.00474650144283328,0.00996819782527925,0.00516786884137543,-0.00221889658023222,0.00207905575097223,-0.0005917159613259,0.00952804655642714
"890",-0.0275349222793877,-0.0312410883207465,-0.0250263109382226,-0.0298694853229787,0.00488450620659098,0.00577083409967027,-0.0307255024186814,-0.022228595179874,-0.013194662610302,-0.0125843292251807
"891",0.00590698585437011,0.00586352739914209,0.00320873996857629,0.0131956991007267,-0.00615021494194301,-0.00260830019048852,0.0114700922044628,0.0142465644207237,-0.00805686994183386,-0.000910226211123244
"892",0.0110912399712348,0.00204003864866631,0.00639630118405954,0.0234932015014728,0.00149712000106894,0.00104592838489515,0.0171137112051383,0.014046865577378,0.00794952887022737,0.00820039019244789
"893",-0.0129975975085294,-0.0171612232159195,-0.0180084068010308,-0.0102296893561314,0.0169440101245135,0.00637363349297915,-0.019258367944358,-0.0132626013683899,-0.00685815676196899,-0.00271126125667331
"894",0.0223215922644679,0.0361053390073698,0.0183386567927388,0.0302494303623597,-0.0115653368313916,-0.00550239359149785,0.0359652571433478,0.0280762165864759,0.00871819609353808,0.0199366670670988
"895",0.00867934869830234,0.0131393565202409,0.0148309993871276,0.00685092276454657,-0.0106100018801785,-0.00323639510596641,0.0117719951325419,0.0136546845894936,-0.00658912368142117,-0.00310973207646137
"896",0.0104154116398869,0.00733009808816965,0.00104370803522813,0.0068044557174638,-0.00170361251024909,-0.000314117404936809,0.0258333346372728,0.00917179908856358,-0.00490997518855973,-0.000891345105075714
"897",-0.0000896160360005505,0.00643727197095423,-0.00521376791936368,-0.00168928461433548,-0.00963692518160064,-0.00345677390003685,-0.000192662175265035,0.00198836918347056,-0.0173995416568441,-0.0107046737841719
"898",-0.00645457034603991,-0.00834293512832751,0.0115303635085287,-0.005560972748342,0.00324295891060555,0.00430904138164556,-0.00153821031307677,-0.00935426079096624,0.00237861858199961,0.00405774690872085
"899",-0.00487227247869848,0.00224356917164492,0.00621757879893137,0.00170196284496682,-0.000302984139184836,0.00209449193695721,-0.00885776576776909,0.00457839958256878,0.0044823519465842,0.0143690478374703
"900",-0.000181538850357321,-0.00167894706013272,-0.00823919939453932,0.00485423840646981,0.0155651725472492,0.00585008669070741,0.00349738132959798,0.00113888918401206,0.0104995799238814,0.0132802587701601
"901",0.0225810754530933,0.0369957360861595,0.0218071667400843,0.0258455454518951,-0.0140381344198846,-0.00309338478504195,0.0303967703223789,0.0301567191024901,0.000432963900475647,0.0192223290506586
"902",-0.00478896510886351,0.00135107236552923,-0.00406529244650511,-0.00470922398077223,0.00577195335990188,0.00470068227307352,-0.00526141200812136,-0.00856107624246605,0.00389472906443888,0.00342901439923127
"903",0.00668352940650507,0.000809791919815783,-0.00204064581456431,0.00141920845710164,-0.0076519038449463,-0.00415811009554823,0.00321117299405582,0.00334259356050537,0.00629367197678543,0.00854337299574337
"904",-0.00106244439195435,-0.000269332519901244,-0.00102248379452896,-0.00448816693291654,0.00466753583598067,0.00480165626405538,-0.0124270032638332,-0.000277637543416476,0.00222757023451359,-0.00465902280095076
"905",-0.00407622942012864,0.000539593520220372,0.00921213106320007,-0.00142402217318394,0.0109065908549077,0.00654566520661581,-0.0032409523825242,-0.000555332933078634,0.0073516240207312,-0.00893604810459558
"906",0.00533873819670272,0.000808562304690064,0.00101415794647508,0.00522813341185557,-0.00369594833999087,-0.000206484488215919,0.00994650610218772,0.00611268318971403,-0.00373382565287939,0.00343490326253937
"907",-0.00539885850008581,-0.00673480388665426,-0.00607922582833265,-0.0137117169304899,0.00210515248465448,0.00505868834704715,-0.00776551668171965,-0.0107707139157438,0.00281091136608325,-0.0106975486074448
"908",-0.027406949878642,-0.0461078766763443,-0.0336391344624051,-0.0318790498483933,0.0134076057268024,0.00564986493934394,-0.0240502745082748,-0.0337797383568538,-0.00331272394514415,-0.0224913537169457
"909",-0.00613022988384337,-0.0025591610839677,-0.00316449176848399,0.00173290271250992,-0.00246806075490358,-0.00255407141421626,-0.0115393415488049,-0.00115589388074067,0.0121868165054311,-0.00752215774694576
"910",-0.00294589240628895,-0.00427581063121185,-0.00105852877239876,0.00543734550125019,0.0124721107061911,0.00430193445002014,-0.0021764069708623,0.000868049107810576,-0.00025258062438116,-0.000891650799776267
"911",-0.000461143416659371,0.006011825259151,0.00741579303736439,0.00934144250607916,0.0250264422993924,0.00723949283832703,0.000991423256227364,0.00289021862725303,0.00833758646349314,-0.00312356292659821
"912",0.0122850477430971,0.0108141275230369,0.00525738098908923,0.0104725137357016,-0.00572227004171222,-0.00506171003864209,0.0217909091400135,0.0193081285599241,0.000167017451757623,0.0143241167204717
"913",0.00182529546295274,-0.000844747131048207,0.00627623457270077,-0.000722885644311777,0.00268608841018092,-0.00101816168577662,0.00019388616940752,0.00452373802366091,0.00392485177453028,-0.0039717927589521
"914",-0.0173969791179439,-0.0166243688050208,-0.00207894891135552,-0.00771855290293599,0.0155935222087,0.00448180434789158,-0.0226787743545706,-0.0115395884260828,0.00141405754937574,-0.0101905157808873
"915",-0.00324445841074006,-0.0160458833102655,-0.00937489638406663,-0.00291667832036757,-0.00113072058257568,-0.00324469701649266,-0.00297500243140836,-0.00740306845909167,-0.00348864526529324,-0.00626679242697858
"916",-0.00381290113938371,0,-0.00630935373299968,-0.00902017901477237,0.000188786005203667,0.0013227179106492,-0.00477427030510569,0.00143408221251784,-0.00158374592328292,-0.00675680343109109
"917",-0.0148430090788431,-0.017181134892331,-0.00105852877239876,-0.0127917022160695,0.0160286608510158,0.00792440037501096,-0.0043975314190644,-0.00887977982523513,0.00484222745735696,-0.0113379006567939
"918",0.00388497787476849,-0.00088897135024868,-0.00317740741390315,-0.0064792588314041,-0.00324790229755201,-0.00453578843375047,0.0130495680550977,0.00780320919670996,0.00830840803997668,0.00504599179799725
"919",-0.00670201103780454,0.000296796213660189,-0.001062811279256,-0.00627040256392808,0.00940296850111566,0.00455645555214268,-0.00554888172797363,-0.00286744222113888,-0.00329599535847069,0.0114102993379197
"920",0.0154901259107578,0.0195670455937351,0.0127659091508847,0.0219587278280229,-0.028315690108109,-0.0114904732736011,0.015942837487662,0.0192692059712718,0.000413384593364707,0.0171480117157852
"921",-0.0145050165729698,-0.0171561926557878,-0.00315131762499032,-0.0165470909200733,0.0191739414346663,0.00764743820324032,-0.00921964392724595,-0.00846504731285447,-0.000826361444072998,-0.0017746899064317
"922",0,0.0056213285570943,-0.0115912057686592,0.00602687876587704,0.0110835401984286,0.00445219575113009,0.0093054367405816,0.00825292322300863,0.00967660211143473,-0.0133332888102071
"923",0.029911563485568,0.0385407357049916,0.027718713900601,0.0351971097178938,-0.0206765997961945,-0.00720083216577083,0.0315806232597584,0.0273776415682345,-0.00319462642210622,0.0198197805590823
"924",0.00931239248794435,0.00821529907113039,-0.00311205922951452,0.00168797957587818,-0.0105661401404264,-0.00417136209428326,0.012550100795506,0.00576957047169646,0.0049305529635868,0.00706713234755285
"925",0.0129717901868485,0.00983397307762957,0.00728378633741444,0.0117956510395381,-0.0123950415705241,-0.00572027822472243,0.0131450931459809,0.0106523675268919,-0.00351623187900707,0.00526322156738601
"926",-0.011272473466112,-0.0178072152762699,0,-0.0145131691803174,0.0204676882182129,0.00791124386920927,-0.0139012792782699,-0.0132429304373244,0.00689312319962965,0.00523562019718837
"927",0.00702306073261383,0.007365361892818,0.00206639461837632,0.0108642392553024,-0.00794731594718345,-0.00275245931303048,0.000563566716175856,0.00520374581880034,0.0000815158944136307,0.00217010912772109
"928",0.0046189360396367,0.00899884432611797,0.00309271934553856,0.00573200284740794,-0.0197409121263471,-0.00787051329051014,-0.00751396557121786,0.00844724768679628,-0.00937169757453915,-0.00563024417114466
"929",0.00504866150198491,0.00641028753881723,0.00719395601643402,0.00356205483580196,-0.00457223940066298,-0.00288502769943644,0.003974451894869,0.00162098381313269,0.00139852749915326,0.0104531334813114
"930",0.0111228962655501,0.016062000517312,0.0102045378083124,0.0238997212064158,0.0048865457069962,0.00475308273773623,0.0156490433777776,0.0148369367728307,-0.000903639179241633,0.00732757416011309
"931",-0.000620716209298822,0.00953950231126832,0.00303032819113835,-0.000462193149210033,0.00962867155089508,0.00503867871314201,-0.00297051973409834,0.00053128995772056,0.0197335466271942,0.00299525195401307
"932",0.00381707808499643,0.000539959362641174,-0.00201448718816566,0.00138733382164635,-0.0148350940938932,-0.00347842289940259,0.00782001360378404,0.00106302975464634,-0.000645016948355503,-0.00170654908078371
"933",-0.000265449640192039,-0.00215867185548591,-0.0131179801687248,-0.00507973960883223,-0.00987554300253624,-0.00349191228669343,-0.00535768717890373,-0.00371550209122462,0.00556716950835612,-0.00512813520556832
"934",0.000373505486599202,-0.0102758735525861,-0.0030675407980153,-0.00162440515485995,0.00404870125993662,0.00226728263595155,0.00297217606965239,-0.00583103961207132,-0.000722105449460941,0.00343637901994409
"935",0.0152901977391731,0.0193989280232596,0.0174359484286253,0.0158065413526796,0.00580299438445797,0.00308440746713878,0.0224071207616445,0.0172975443636474,0.00264976712180998,0.00813358273024756
"936",-0.00201351447387788,0.0026802593837294,-0.0110886775977176,-0.00297514222772555,0.0138862961529582,0.00932703272033408,-0.0157578630374883,0.00239127540918616,0.00912948644679701,-0.0106157845556669
"937",-0.00491338639108108,0.000267415330798437,-0.00305813014536649,0.000688797238427741,0.00896991487624588,0.0015227358193175,-0.0103056211421821,0,0.00150777713661165,0.00600867863313748
"938",-0.00811172576270114,-0.011758507982219,-0.00408999478773486,-0.00642195338898288,0.00286760841488132,0.00141955212861711,-0.0224321805476352,-0.0108667748853657,0.000792440589360677,0.000853142814789987
"939",0.0206225455714357,0.03163890952696,0.0133472670440409,0.0184672062548359,-0.0134395480778881,-0.00496062661354901,0.0272446500089869,0.0262591161867489,0.00308787799474564,0.0153453669436308
"940",-0.00479003238304565,-0.00655317907483377,0.00506562282775347,-0.00181321026638681,0.0173908489597736,0.00773257635917912,-0.0098988659922975,-0.00626607060462714,0.000236790587468727,-0.00671712532960733
"941",0.00350048585500096,0.00897101811986567,0.00403239064876781,0.00726618264917667,0.00683751755562079,0.003331875612955,0.00264097728867463,0.0105095742037511,0.00891727423518573,0
"942",-0.00174410062842478,-0.0047072037787419,0.0050202008238367,0.00338138215219974,-0.00415007030346826,-0.00241532768290453,-0.00733801598931549,0.00052017906575097,0.000782158792055565,0.0131023214391592
"943",-0.00297018093883061,-0.00551769917028855,-0.0119880828243185,0.00584136752952835,-0.0006633908142335,-0.00121044681857052,0.00227460008400304,0.000259663758453321,-0.000312567416472787,0.00584064025226727
"944",0.00420539798179753,0.0105681523103975,0.00202198661393216,0.0147418683601708,-0.0048319726734527,0.000536800766123058,0.00491690835184455,0.0161084250254995,0.00781799678467676,0.00207379995796053
"945",-0.0075036475293766,-0.0138563431980826,-0.0191724348168922,-0.00308149840497129,0.00258109702722331,0.00354141118658813,0.00846816037853282,-0.00946088768658759,-0.0034907841597771,-0.00331121313906824
"946",0.0201317249763939,0.0291624239664614,0.0318930467844596,0.0181054265873093,-0.00600723664339275,0.000201551975886671,0.0130618923317167,0.0216833115846053,0.0196948300026172,0.0203488153415423
"947",-0.0000860836387882591,0.00566714026010628,0.0109672985443989,-0.000433752386613806,0.0125657819675005,0.00645167582907602,-0.00294674147112561,0.00757941396955775,0.00625996617070146,0.000406994849060593
"948",-0.001206527386443,-0.00179297359243713,0.0039446717968501,-0.00889555674455345,-0.00833661649561412,0.00100175382516365,0.00221652836472774,0.000752248485863083,-0.0109248389488635,-0.0101708574073451
"949",0.00560883406520207,0.00487543243043231,0.00491147994297214,0.0120404332777733,-0.00439346824753473,0.000399941422157379,0.00129031962110493,0.00651448572636193,0.00989498388797205,0.0332921999423756
"950",0.000943699046664248,-0.00229840928491554,-0.00195498438386033,-0.000649561821143396,0.000190901144288658,0.00100054527018956,-0.00147235949163049,-0.00174237527229026,0.00478496871380951,-0.00477328649540332
"951",0.00308627329317268,0.000256087249669301,-0.00881490492568404,-0.00411210544642204,-0.00988086350075823,-0.00289814190602466,0.00866487087903733,0.00324195951788564,-0.00249441391987992,0.00479618003680238
"952",0.00777699289318301,0.0174000511435404,0.00296425041358894,0.0184742624928946,-0.00154967138488915,0,0.00987027240883176,0.00870020622403844,0.0159896929984249,0.00477332743478698
"953",-0.0039005672692366,0.006036180565266,0.00689670719924051,-0.00170726652359032,-0.0149443970669204,-0.00571181075777227,-0.00307671964848988,0.00689971701152658,0.00507192484893348,-0.00158359108553852
"954",0.00204300995877649,-0.00249961638537677,-0.00782758905414171,-0.00128238457380958,-0.0122155897351429,-0.00433383894298867,-0.000544905709370491,-0.00587373404045455,-0.0079406827458256,-0.0111022708620921
"955",0.00492783548100806,0.00375944874077772,0.0069031900178087,0.000427984198095199,0.00807855025390758,0.00475787688416585,-0.00508593536573476,0.00787791818347494,0.00448837545944514,0.0100240858846563
"956",-0.0131042282131049,-0.0269664138938888,-0.00881490492568404,-0.0316647719630234,0.00603427391380285,0.00342550263152441,0.00492953218929104,-0.0315094278424444,-0.0310544982950141,-0.0293767432883081
"957",0.0097658666785263,0.0197587111434996,0.00790505181569512,0.0159080206399234,0.0021638887561084,-0.000602751174311078,0.0199855105905735,0.0214372659555819,0.0092998692698496,0.0237218936144195
"958",0.0022054803301701,-0.000503140776916045,-0.0127452168321784,0,-0.0118735867316322,-0.00552551438659521,-0.00195962599778643,-0.00864169694159933,-0.0140877695810663,-0.0123852560833844
"959",0.00186269200500888,0.00075502461905308,0.00794441974505511,0.00108756686278655,0.00675276399142821,0.000303330855733197,0.000178504568216109,0.00498120715874584,0.00200814859034404,0.0084953217711945
"960",0.00295745560751381,0.00327052252051452,0.000985182346324942,0.0108626301737067,0.00286085024746718,-0.000303238874026168,0.00196309772374925,0.00272631493914433,0.00863339269662822,0.00521452919396115
"961",0.000168237614001754,-0.00802404426394199,-0.00984238538390314,-0.000859542681096448,-0.0154422840090231,-0.00666730162211027,-0.00587711777414734,0,0.000229262503816718,0.00518756107376728
"962",-0.00286347612899962,-0.00910017759455184,-0.00298204597787133,-0.0169931590021656,-0.00879094863775143,-0.00579642097993049,-0.0100326047676567,-0.00543742209540188,-0.0103912052876222,-0.00317590168457615
"963",0.000168774216145584,0.0104594023990416,0.00299096517353714,0.00634584909722125,0.00272101023537186,0.00583021536257555,-0.0061524562577685,0.00447298225618287,0.0132798096578193,0.0051772725314605
"964",0.000759657601346442,0.000252529308628846,-0.00397604198699419,0.00282678678649595,0.00934783372998793,0.00447476769864341,0.000728371211032419,-0.000742198574226416,0.010515010266877,-0.00237718728795866
"965",0.000337930408804477,-0.00631010632471185,-0.00998016319365225,0.0110582992357275,-0.00430599881673566,-0.00167400582764377,0.00727763003142678,0.00396151703237702,-0.00527821615435886,0.0063542032704953
"966",0.00793057830068822,0.0182879883078753,0.00705652202236839,0.012438042045555,0.0131428899426433,0.00335446178806365,0.00559996827447629,0.0133168274917279,0.00432085361311185,0.0090765567807225
"967",0.00401766113051294,0.00698435139687681,0.00300305776704235,0.00614277444203215,-0.0203998971872447,0.00324199515486301,-0.00107795333149063,0.00219020568116446,-0.00694390493833852,0.00469301607448758
"968",0.0192580994493996,0.0240277576284647,0.0229539855270935,0.0227369757956686,0.00778447520152836,0.00807878425262865,0.025894888367451,0.0182126060604542,0.0338982424771019,0.0237446438397573
"969",0.00376241056141158,-0.0128206045153749,0.00878050617176118,-0.00185253040570332,-0.0171531444230943,-0.00420768816365047,0.00999133964064214,-0.00310009791207866,0.00257300597348387,0.00418253064980045
"970",-0.00187411446413677,-0.00833120158548339,0,-0.00412482915765822,0.00449069044985317,0.00030229804559978,-0.00485956005961785,-0.00956969517930262,0.0102653904434158,0.00265047491442716
"971",-0.00718433075205871,-0.010377910529408,-0.00676978044298193,-0.0126320539538284,-0.0220482153384604,-0.00844790685737307,-0.0361003784152456,-0.0164250098592188,-0.0158949268100952,-0.00679756808052623
"972",0.00402903276480782,0.00124808255082787,0.0116845606292368,0.00734058155227002,0.0013507101660839,0.00375227659796673,0.0119411781769598,0.00171905200550504,0.01216910575025,0.0106463598290467
"973",-0.00376734197183504,-0.00997484760503198,-0.00577486037398656,-0.00978546707123573,-0.000518803157333547,-0.00111167576987958,-0.0080455333845334,-0.0132385608982362,0.00306032486664498,-0.00827682583247247
"974",-0.0118382854908138,-0.00554175374992771,-0.00774446220667913,-0.0241797679262798,-0.00539821906180615,-0.00829573525020466,-0.0093727852422385,-0.0134160862352553,-0.0288391826575858,-0.0417299075536764
"975",-0.00141406417402856,-0.00202598450419589,0,-0.000431238585529958,-0.0208748185873855,-0.0128526017025825,-0.0109171476717946,0,-0.00949961837834368,0.00158342810595902
"976",-0.0155796386766255,-0.0253809586058716,-0.0175610976579705,-0.0262990386988423,0.0248379681386421,0.00744076851621811,-0.0314566515087366,-0.0198944596080615,-0.0109499850619239,-0.0296441914335533
"977",0.000508044677999253,0.00364574750559443,0.0148959172811451,0.00509243320727371,-0.00551331001331978,-0.00287234791606628,0.00873649894984618,0.00179895405660058,-0.00450481786283241,-0.00773932753243955
"978",0.014718099284948,0.0238715205682025,0.0254402633801007,0.0237882775835598,0.00407912043299308,-0.00236619238256597,0.00696661069705184,0.0159013191521238,0.0131154389816137,0.0270935643193935
"979",0.00275089931926575,0.00380133533778726,0.000954188096101705,0.00064556784609171,0.00614586842365727,0.00206206291903022,0.00467454253437105,-0.00530184983282889,0.00083277313446195,-0.0143884167031987
"980",-0.000830995843903115,-0.0143904049792994,-0.00285969652977014,-0.00301012732086914,0.00424460241509306,0.00535108514760707,0.00204741731838309,-0.00380693402284982,0.00968229220156491,0.00324407562208728
"981",-0.0144770794993561,-0.0330428161620526,-0.0191204429592833,-0.0317015256288428,0.00494914528656287,0.00204658185508455,-0.00705802440718351,-0.0236941359342774,0.00696739607334118,-0.00242518921933998
"982",0.0147737694556116,0.0105959340503494,0.0175436657604213,0.0231622193676602,-0.0178505856716022,-0.0107250872736823,0.0192671192631304,0.0120041452142881,-0.00171126399192723,0.0186385273102563
"983",-0.0116470571116382,-0.0152030765155502,-0.0162834597294108,-0.0248146905786233,0.0138922184268795,0.00433700932945325,-0.00293621351348006,-0.0128933507888794,-0.00797430359084894,0.00477332743478698
"984",0.00303026561527941,-0.0167690197739486,0.00486863788576541,0.00781269425174647,0.00855014146892485,0.00215894148770412,-0.000552401511870193,0.00261236111693375,0.00300498833292018,0.00197938699468603
"985",-0.00562297167664993,-0.0151596843935038,-0.00484504909617733,-0.00819518551117593,0.00520950151073962,0.0017435316997767,-0.00386736742924787,-0.0122456757579326,0.0143060674970439,-0.00948249177806404
"986",0.0212680363762283,0.0321605366586462,0.0204478533787145,0.0285843520282469,-0.0222296921303963,-0.0131499434816271,0.00758014809996554,0.026905431622031,-0.000295325657883816,0.0295174429557872
"987",0.0128085946249683,0.022902870610759,0.00954199221713381,0.0197567175372309,-0.00260677314928737,-0.0024968499268565,0.0135776976708275,0.0215773052748895,-0.00132964982531958,0.00852383101731813
"988",0.00269292703727642,0.0119758980969942,0.00567104333923307,0.00361929880235912,-0.00784218909790013,0.000104932858573825,0.00144812256454108,0.00578321809282456,0.0212278850864176,0.0126777038589156
"989",-0.00105810755335611,-0.0100335274974481,0.00469925193099119,-0.00169704811419891,0.0141220458931499,0.00625570258552544,0.000542335031401997,-0.00399984089391814,0.00753236725772033,-0.00113815050425914
"990",0.000570299828820175,0.00571766128673734,-0.0121609296649855,-0.00467475067333123,-0.0214063659592751,-0.0165797618129927,0.00325203966302845,0.000251015579069813,-0.018762137741628,-0.0068363323991949
"991",0.00366362625227667,0.00594290655403618,0.0028408231442123,-0.00640493727427993,-0.00966391842611425,-0.00853557448902797,-0.0149468882529212,0.00250952586061226,-0.0125275238095237,0.00764819747851098
"992",0.00389372054208392,0.00154154036789533,0.00188874652894411,-0.00343782707088336,0.00493269352631032,0.00212576340660964,-0.0107860135773189,-0.00150220467588225,0.00430300489740354,-0.00265651027620528
"993",0.00581763871156249,0.00461581034122971,-0.0028275453134603,0.00452795270883555,-0.00608207185877319,-0.00848465817541388,0.0103494747750981,0.00350951208472372,0.000295552939925781,-0.00152208837496137
"994",0.000642666586721408,0.0104678218261363,0.0132325079279085,0.00643909533651832,0.00375712245333393,0.00320936105457714,0.00256068195694881,0.00949289118139363,0.00472637900520279,0.00990851900668721
"995",0.00088316101024577,0.0015158574078884,0.00373157461278462,0.00149278819853871,-0.0145453638852763,-0.0105561714163451,-0.010217297092379,0.00445450708381179,0.000955457531301773,-0.0026414734242225
"996",-0.00457206079692773,-0.0151362632980371,-0.00650582903361585,-0.0161844034804673,-0.0130231973948143,-0.00409429426714147,-0.0110595284394954,-0.0101010957102814,-0.010867940050489,-0.00264846928545504
"997",0.00580169031702416,0.00512297489583391,0.00561298846971603,0.00281423052749119,0.00692725460094845,0.00595069387400415,0.00260925914443,0,-0.00660726815012469,-0.00341429533432092
"998",0.0010711498500533,-0.00713554203037303,-0.00279093780369288,0.00151133400100978,0.0182377990248523,0.00860503600258644,0.00780804402826951,-0.00971614631604945,0.00291457294543851,0.00761322130876096
"999",0.0024134044654176,0.00268691930355369,0.000932825674877957,-0.00452631575615015,-0.0010729551052725,-0.000106417341430243,0.0114371848562906,0.00510720690557753,0.00678095395188438,0.00906686105773313
"1000",0.00634017151135846,0.00541073021610949,0.0059117804158122,0.014597219347591,0.00697890680663393,0.0021332577513915,0.0109428497146409,0.00909325583847886,0.00155433349452783,0.00636464767940859
"1001",0.00311038387557616,0.00358805484638447,0.00373119464799343,0.00344073570503589,-0.00714337096278372,-0.00276741896971566,0.0069659739293253,0.00715624251854252,-0.00199529992634417,0.00520837720647793
"1002",-0.0014312438618177,0,-0.000929277334719147,-0.00107153487707412,-0.00204080800982775,-0.00352177426246369,-0.00307874774137362,0.00131573857957457,-0.00288781185736087,0.00370098782268258
"1003",0.000398377934979433,-0.00689484572483401,0.00279045201390704,-0.0032182874105976,0.0089318902791462,0.00385573232454317,0.00799269393923763,0.00630759305385009,0.0026733995938395,-0.0018437084596814
"1004",0.00143264777577845,-0.00128583277187244,0.00742109860909435,0.00086112725688392,-0.019584729359627,-0.0105050773128568,0.00396501565670571,-0.000522166564960513,0.0162938596861544,0.0107130102608699
"1005",0.000715150693035183,0.00926878107851081,0.00920840604244177,0.0128025176148043,0.0169195696015922,0.0112433250222188,0.00448737508901575,0.00966804867489368,0.00357095173028021,0.00036549207135006
"1006",-0.00158842826563699,-0.00459176296734809,-0.00821195970789912,0.0050989197445217,-0.000751745232832168,-0.00203121289341213,0.00125083074337629,0.000776342423359333,-0.00493797084768133,-0.0120569444895691
"1007",0.000238662475757989,0.00666336239226251,0.00368002706406712,0.00697498554383214,0.011064397667252,0.00503449391383115,-0.00124926812040449,0.00672391330356992,0.0123330804373718,0.0188608017722003
"1008",0.0103381867836703,0.00814684838775515,0.0091659903300112,0.00965589853641835,-0.00754365231200071,-0.00309079253084643,0.0155468230785389,0.00899010298037473,-0.00519031859003516,0.00435584443840731
"1009",-0.000551062029188754,-0.00202031962901017,0.000908281692594048,0.00457374518988152,0.0011779838250694,0.00235263609795755,-0.0177721835715844,-0.00509132980444837,-0.0235507246376812,-0.0133719597444494
"1010",0.00519745784144865,-0.00632607670756646,-0.00725947582680109,-0.00248318094164723,-0.0220274581762469,-0.0107732523459172,0.00412015438893265,-0.00230325696904654,-0.00282007421150288,0.0106226410499182
"1011",-0.00195845883998547,-0.0114590439517531,0,-0.0105809301581744,0.00437339807845083,0.00517530998254556,-0.00535227273358396,-0.0143626286573442,-0.00401870224077916,-0.013410585848192
"1012",-0.0019625194713534,-0.0054092019670513,0.00365597626670588,-0.00922610591624673,0.00533447701468903,0.00665067724272062,-0.000358802544160541,-0.00312267378608166,-0.00186804151732733,-0.00367371914114689
"1013",-0.00125837838940257,-0.00492151551009479,0,-0.0103708640254304,0.00541394036993492,0.00341054773041316,-0.000358652045159502,-0.00313232949297204,0.00404246887194981,0.0117994381284996
"1014",0.0035438821366407,0.00702757884305316,0.00728602949005097,0.010692864315774,-0.00560009305480191,-0.0039292126713294,-0.0017953259349901,0.00418966066683546,0.00589031486319391,0.0112973335278741
"1015",0.00902457192474526,0.0294651696818202,0.00904178340455131,0.0201018283725107,-0.00779809370705475,-0.00287943698013093,0.00449600565392427,0.015124212498125,0.00407681405153615,0.0064864718915163
"1016",-0.00163321473317768,0.00477047390941499,-0.000896384918070869,-0.00871203283485567,0.00895059335263171,0.00673645822292213,0.0028641592337979,0.00154087017485138,-0.0104090058108441,-0.00143220592840976
"1017",0.00724447120517935,0.00924517375447276,0,0.0029297109414359,-0.00638332007461617,-0.00276097046826085,0.0067831780518377,0.00641177584430319,-0.0101454753417649,0.004661289919627
"1018",0.00170154043019455,0.00990350005443164,0.00269084041909529,-0.00146052575026678,-0.00468134442877244,-0.00244980678120088,0.00939711834047463,0,0.00557684067259268,-0.00107079602915094
"1019",-0.00980544970350838,-0.00833556501093868,-0.00178883779715866,-0.0077310793926656,0.00721951344995708,0.00256160806551153,-0.0119442675575983,-0.00535150809844731,0.00217348433796283,-0.00107179677897651
"1020",-0.0013256160528573,-0.0064277970947878,-0.00896076213419417,-0.01094964900665,-0.0137939296884676,-0.00777312592882073,-0.00213342719084797,-0.0102486648854151,-0.0188453782617007,-0.0100142801895847
"1021",0.00226444463405739,0.0126898027904305,-0.00994546178101163,-0.0104319940950391,0.00792971010936694,0.00332667596867897,0.00391950261291774,-0.000258598062970572,-0.00129571649304228,0.0101155804464559
"1022",0.00568657480806345,0.0100739090784427,0.00639262442895894,0.00774541238028026,0.000436868999990958,0.000107147347286451,0.00496869430806091,0.00699082426468789,-0.00511331759988787,-0.00858361088916537
"1023",0.000542162388881939,-0.00267586023247635,0.00907449584251441,-0.00597794857861222,0.00950214186161413,0.00502714754413702,0.0105951106458497,0.00539987740407599,-0.00199443846276126,-0.0126262752838782
"1024",0.00387101642853449,0.0053657275153578,-0.00179880188006187,0.00880564976571074,-0.0151464316543403,-0.00606622118986178,0.00279594273566297,0.00332486088319128,0.00814756303700692,0.0222871715082313
"1025",0.00246780060546503,0.00558011463477004,0.000900839126991348,-0.00340625887598467,0.00450403824432022,0.00374737881670262,0.0139397992842674,-0.0025491760771218,-0.0246264402370709,-0.00857762194444589
"1026",-0.0174630035545229,-0.0243669366092848,-0.0171014766781417,-0.0316172581419635,0.00524918004158037,0.00458758638761925,-0.015638392495766,-0.0171222706644715,0.0183694129602125,0.0126171730460689
"1027",0.0075164928293856,0.014095160084499,0.000915581915736707,0.0105890713208565,-0.00761496117762361,-0.00392870599930606,0.0118712068616489,0.00832011979199621,-0.00314709858111084,0.0156639803234693
"1028",0.0160085474003779,0.0246281806476947,0.0201278729754708,0.0242304221349945,-0.00495081408050446,-0.00465011833233497,0.00465849362328341,0.0180510084404768,0.00716106903677027,0.00736068056253858
"1029",-0.00191188322456026,-0.0033317614925642,0.00986567919949755,-0.00745959369500482,0.00022164618149545,-0.00236204236548954,0.000171578369860148,-0.00303950129710662,-0.00267588678877939,0.00974249329415966
"1030",0.00222219753739683,-0.00501469328836901,0.00799288705249346,-0.00128831202737967,-0.00829077649538623,-0.00570472197994742,0.00257554208771293,0.0015239550203654,0.0134151018799946,-0.00654715488960811
"1031",0.00282923291739245,-0.00287941927856117,0,-0.000215039152968499,-0.0101430419133369,-0.00616999391424811,-0.00907704855468316,-0.00608817624282987,-0.00408466726364609,-0.0055498412586894
"1032",0.00625203974367672,0.00601672062435687,-0.000881175411374779,0.00129051242851119,0.00518063078696063,-0.000435723557833056,0.0112342599785713,0.00280756143282468,0.000151822872495266,-0.00279037104622348
"1033",0.00454676393725295,0.00717680187881919,0.00617315736797641,0.000429668528459271,-0.0091854117521849,-0.00686447664598522,0.0025634875057341,0.000763662750517646,0.0110875309660747,0.00664576963206298
"1034",-0.00226291498991749,0.00190044244500465,-0.00701164722392533,-0.022971425658562,0.00870435592999264,0.00570557029268559,0.00238680513336531,-0.00940979331279668,-0.000525702272237361,0.00486435090443704
"1035",0.000378079255538122,-0.0101943674070495,-0.000882322098005983,-0.00944818158633942,-0.0115438320274305,-0.00327318770759955,0.00323132313707841,-0.00744582215201461,-0.00165327262664072,-0.00587820501003333
"1036",0.00597026360906705,-0.00047899922895267,0.000883101277778131,0.0122003568346942,0.0144007336762526,0.00459725640430131,0.00627236685117549,0.000258896585580759,-0.00398945409155649,-0.00347824910264893
"1037",0.00240395242757274,0.000239582964746132,0.0088264150218289,-0.00504051247923776,0.000669789379646568,0.00032649717849309,-0.000168478983748388,0.00206872366037936,0.00476110917980832,0.00488653099623337
"1038",-0.00314762760315646,-0.00167727597839318,-0.00699935282454933,0.0019823224156581,0.00446911345035317,0.00228757155983117,-0.00336990906514367,-0.00567747366345184,0.00767208742396597,-0.0128516878535987
"1039",0.00631547712676639,0.0112794484953975,0.0140968935340076,0.00835343075898143,-0.00322524258635681,-0.00141287930666989,0.00287402446336782,0.012457736235713,0.000970403814507748,0.00738913410732644
"1040",0.00298816492356524,0.00427140612878651,0.00868818093788182,0.00348804907457079,0.00156181346555306,0.00370064101735057,0.00134876472519752,0.0084595133516665,0.00700959700180781,0.00314354882990564
"1041",0.00208574485315971,0.00472609634698329,-0.000861342143217869,0.00608311907359504,-0.00311854182941873,-0.000217162377157631,0.00387193062540048,0.00279630606525805,0.00274001050933093,-0.0010444823480118
"1042",-0.0200699083696808,-0.0275166875115673,-0.0275862859001982,-0.0319585174044522,0.0149727967928961,0.00965155032288911,-0.00905574603961046,-0.024081443510435,0.00649870005173336,-0.0013942307795789
"1043",-0.00614419549144096,-0.000967233954767166,0.0017731847993343,0.000892147015820077,0.00363405960898122,-0.00247051798679709,-0.0079542392206009,0.00545478650174558,0.0089515156112745,0.0223385505785685
"1044",-0.000687107123407804,0.00145211275358403,-0.00265501803019341,0.0024515894412025,0.00636222124020747,0.00258412702228883,-0.00545875969207443,0.000258520575192822,-0.00749035733729753,-0.00887669868527741
"1045",0.0106928538143729,0.00991066467220936,0.0133098387489559,0.0120054266285816,0.00588621180956239,0.00322202331502264,0.0178388417742295,0.0178198945684758,0.00659443893887568,0.0220461048357377
"1046",0.00619663624495081,0.0117282483167185,0.00963214573999904,0.00593134308241949,0.00130046213557833,-0.000427476290448592,0.0208965764751476,0.0134485543483476,0.00203813502554451,0.00168514618857385
"1047",-0.0166730457922277,-0.0160870831376146,-0.00173466215041007,-0.0102642738282822,0.00289863866529494,0.00113781440638827,-0.0269065260068795,-0.0160243889888628,0.0172162932669973,0.0151413553204189
"1048",0.00213862413852173,0.00673213432473152,-0.00868787910510804,0.0136803624396857,-0.0153732728873859,-0.00525444439320533,-0.00797303349858358,0.00508943585450239,-0.00078555310137518,0.00397754323492205
"1049",0.0172241947993419,0.0128973253635372,0.00964056138747993,0.0198086385202902,-0.00978506470205065,-0.00679083122113922,0.0143639153913002,0.00860739125352872,-0.0130789167106762,-0.000330205386527171
"1050",-0.00749200419442386,-0.00848870401169954,-0.00694457079699617,0.00106718539264761,0.00832795762073779,0.00716252395808303,-0.00859736435462788,0.000502214697388537,0.00912455671300028,0.00495373116318754
"1051",-0.00785098132491313,-0.00808557879988625,-0.0192305901376388,-0.0140723890068108,-0.00638736140911977,-0.00247798507029773,-0.00646154664927168,-0.00777707179900911,0.00265514879131024,-0.00460062643848858
"1052",0.0087498417313514,-0.000239509233068369,0.00445612498958536,0.0134081999990496,-0.00609544870850187,-0.00237704306146691,0.0124934398125931,0.00227556065744494,-0.00257658171645725,-0.00858377702770841
"1053",-0.0014331947736318,0.000719297335844971,0,0.00192056013271746,0.0097012283314768,0.00584803315058235,0.00050709794818582,0.00327936368433734,0.000358804532442303,0.00399601803386762
"1054",-0.0185056548004114,-0.0230050868642229,-0.0248444569118673,-0.0296059991905143,0.0167862631526821,0.00850445188132998,-0.0155429624902571,-0.0226302164836151,-0.0117638616522814,-0.0162520558719252
"1055",0.00692602851548485,0.00392445841325606,-0.0163784531123174,0.010316091895834,-0.0056477430468771,-0.00234849427499151,0.0113265000184428,0.00102903974742041,0.00326629155066294,-0.00573161612253437
"1056",-0.00603759515596292,-0.00464217084339535,-0.0703056008385818,0.00586573201748442,-0.000436893220821077,0.00224725289482963,-0.00678766206782155,-0.01876127952152,0.00463029948900107,0.00271274688097622
"1057",-0.0114574366680056,-0.0252822809014642,-0.00198985581438405,-0.0166307293620629,0.0149706218526369,0.00362973018673185,-0.00803005384208322,-0.0275010904723966,-0.01865185785214,-0.0365235273160286
"1058",-0.0185127323079621,-0.0307226474717129,-0.0368892224178861,-0.0204259516759282,0.0113056178134379,0.0085093548658941,-0.0130899565818412,-0.0250473026786308,-0.000220143825636065,0.00596703307699742
"1059",0.0132352557526152,0.0350741229331366,0.0455485469612613,0.0123318546760607,-0.00766601247469545,-0.00305871583376482,0.00837716056530202,0.0256907876120009,0.00535816187029647,0.0310536687711132
"1060",0.0036371097057557,0.0107930990023966,0.0267329003384578,0.0017719706167878,0.00268224200509315,-0.000635119730110767,0.00882621265162964,0.023739064794849,0.0102211724449064,0.00575298742614816
"1061",0.0154979274327744,0.0245840816440703,0.0289292297707175,0.019234893627871,-0.00588489820593574,-0.00518693566317741,0.0109797400217626,0.0237972489618687,0.00556481916473284,0.00471070698178733
"1062",-0.00346851551828231,-0.0026658463312822,-0.00374867998493578,0.00303698041679157,0.00333637476512672,0.000532073133469924,-0.00899370266255084,-0.00723154011171878,-0.000646801787025919,0.00736764965761338
"1063",0.00286170791822427,0.000728847527653009,-0.00564453225003458,0.0131919840155588,-0.00128687104927905,-0.00127670150885073,-0.00753432905252416,0.00884473615366854,0.00927718786169329,0.00199472211951734
"1064",0.00956317703937426,0.0150558483343455,0.00189229171322336,0.01152610490883,-0.00751845161958287,-0.00511130629001921,0.00465849362328341,0.0105725184083938,-0.00798058309763683,0.0033178730098975
"1065",0.0030563420265588,-0.00885176440470914,-0.0245515532480585,-0.00105522998698504,-0.00248959288666084,-0.00267623305416265,0.00507559483943965,-0.0109720465798473,0.000287271941622924,0.00264546644963271
"1066",-0.00243762341037301,0.000724175120414339,-0.00193603158814337,-0.00506953130144527,0.00141078168858622,0.000321473457763455,0,-0.00438606376752437,-0.00517019981222888,-0.0135224126400227
"1067",0.00671867242708335,0.00410022549927613,-0.00194001171959379,0.0114647458138388,-0.0076924074688115,-0.00289675177396409,0.00448103641202002,0.00103630290046652,-0.00238188260916128,0.00568367458562014
"1068",0.00690116241179717,0.0100889257470753,0.0155491923207081,0.0128043904902611,0.00797001384685814,0.00344398129877721,0.0116680146843267,0.0111314364055637,0.00332820328993977,-0.00132973490910149
"1069",-0.00135573861441918,-0.00546965991588777,-0.0124402512496353,0.00870481199162931,-0.00205808680649056,-0.00257389599296365,0.00746244474831714,-0.000768264164570986,0.00858154624044927,0.01564586580112
"1070",0.00422365192235175,0.0119561291263703,-0.00193790762195223,0.0160263110170549,0.00486119652824923,0.00213434424579217,0.00235687700053466,0.00922420844538374,-0.00471903328529233,0.006882928416728
"1071",0.000826074781107966,0.0054346079715164,-0.0135925079180407,0.00849347333149941,0.00108497853954059,0.00225929072502806,-0.000839402444597903,-0.000254199790392873,0.00459769406460553,0.00911459275608784
"1072",-0.000149867656515146,0.00258527206394166,-0.0196849178741966,-0.00200504573113747,-0.00400906195932571,-0.00504469615071046,0.00168085190766853,0.000507919394195699,0.0158038262529698,0.00096772869811601
"1073",0.00315228458042593,0.0114863764256454,-0.00903610658100951,0.00542484862919634,-0.015012908612329,-0.00431539148479332,-0.00134282528415375,0.00736046292430115,0.00232313969046527,0.00290047881931033
"1074",-0.00254393953555199,-0.00370793791497726,-0.0081054299279214,-0.000999347410009066,-0.0019882083291678,0.000108599864343306,-0.0104181374242232,-0.0136054199636111,0.000912979318971052,0.00192792795831886
"1075",-0.00345035364570356,0.00790868919902898,0.0194076188436016,0.00100034710429697,-0.00531272806418326,-0.0029246835877903,-0.00747150584889344,0.0107280696577647,0.00806967258682434,0.0237332348437118
"1076",-0.00301063894782472,-0.00138481025039816,-0.00701415624133539,-0.0117906740885143,0.000889959842450105,0.00130415380787241,-0.0010265516535235,-0.00732904189155559,-0.0071001320590246,-0.0184837784171399
"1077",-0.0074739075803425,-0.00970647782941825,0.00201831746969927,-0.0188070380335835,0.0107832986693817,0.00564235249326073,-0.00205497285413037,-0.0078919584794469,-0.00722096191265387,-0.020427623687187
"1078",-0.0000761593752368617,0.000933344517880297,0.00402815428060643,0.00824426054646432,0.00626872703106462,0.00388407647342626,-0.00120143530932393,0.00307912718415015,0.00204782852872087,0.00782006312591998
"1079",0.000760720912424961,0.00349728272958294,0.00702122066997179,0.00306628405921128,-0.000765029741824352,-0.00333230711072907,0.0135741742319899,0.00818630552762989,0.0134602119856329,0.00258645032519977
"1080",0.00364852607802812,-0.00232327437266466,-0.000996034001490065,0.00122267522249064,0.0135624681874917,0.00733294987845245,0.011018580000896,0.00304475000976412,0.00862252289301879,0.00515972166490997
"1081",-0.0112085654680379,-0.0251512101191927,-0.00299099463048014,-0.0250357405294391,0.00226526104399194,0.00246225874127548,-0.00989306036000914,-0.0146720722813081,0.00606680442467833,-0.00609568631687829
"1082",0.00574429420939682,0.00860001718612513,0.00299996751721565,0.0144049494200398,0.00430726320480734,0.00128207479831777,0.00778998617267357,0.00770220137425159,0,0.000322850943261122
"1083",0.0136317905486874,0.0272383005129797,0.0149552040659724,0.0236677305042854,-0.00643268069578573,-0.00394615724305547,0.0115949870406764,0.0168152627572835,0.0039060304758598,0.0158115350310737
"1084",0.0051091607029492,0.00691745350944095,0.00392945790930943,0.00884585807315075,-0.000862949024572401,0.00074949693434756,0.00714296848944507,0.0107743035418315,0.00163825938566542,0.00730619171549063
"1085",-0.00104659184178135,0.00160293787462651,-0.000978576081577809,-0.00817040775376632,0.00377968300089782,0.00353068548983249,0.00494767337748603,0,0.000885852498096806,-0.00283811777633758
"1086",0.00860504507716198,0.00983032902706782,0.000979534630738632,0.00863947437388535,0.00968269138989353,0.00426446238175893,0.00935517685181186,0.00793255796704528,-0.00333621581453702,-0.000316316289468599
"1087",0.00652896565366445,0.0178856627576578,0.00195667059437943,-0.0017927054119149,-0.0102289586199876,-0.00286611836410811,0.00455288717006708,0.0108213911863557,0.0192648715922641,0.0060107715714699
"1088",0.00324290503877744,0.00400361008587491,0.0263669882965585,-0.0081818209126433,0.00764328990671825,0.00383298842614033,0.0111686738652641,0.00389295633359565,0.00415556308623799,-0.00723270247891861
"1089",0.00235114607110876,0.00443038108906135,0.00190287435120684,0.00603607724150623,0.00309815929946056,0.00201493167459343,-0.00480252841518813,0.00484721835024793,0.0170203436180589,0.0104529163490235
"1090",-0.00153935506636504,-0.00220541969482124,0.00284916538259927,0.000199956541742541,0.00160493190067057,-0.000307530866120564,-0.000160534902747145,0.0014469270157631,-0.0128633659140043,-0.010031372377705
"1091",-0.00359708428608074,-0.00773652289907767,0,-0.0221955693769957,0.00565961353151256,0.00265354950884955,-0.00675668219580672,-0.0093927278402598,-0.00352369513932049,-0.0104496070956075
"1092",-0.00663082724301078,-0.00757418407291444,-0.00189375470261888,-0.0165642693427077,0.0044598952831798,0.00254183027446397,-0.00550708202218952,-0.0111840809227076,-0.0143448687501713,-0.0160000118565692
"1093",-0.00904828813644121,-0.0255891275496397,-0.007590297684687,-0.00956546441779804,0.00951454034735444,0.00496315714888551,-0.00146613114822414,-0.0118025061751489,-0.0288363576480433,-0.0669918253132131
"1094",0.00441583939396994,-0.00483740588071691,0.00573646387162552,0.0130167003533308,-0.00439843139702423,0.000526024510200784,-0.0053820753692807,0.00870859123509948,0.0127552937007369,-0.00313697441194594
"1095",0.00387487007712584,0.00555512045980122,0.00380193679636798,0.00186533302894398,-0.00105140002276682,0.00146965416971567,0.00393568292712332,0.00419340604866525,0.0143152233795893,0.036713179193959
"1096",0.00853619438784303,0.0112804943026223,0.00473485282044739,0.0117915040198919,-0.00715946235822695,-0.00482413533578496,0.013884293241043,0.00245643184056044,0.00352821944876425,0.00910628911108069
"1097",-0.0105249301704181,-0.0168454453168558,-0.0169648643793158,-0.0220812214174856,0.00572639603359293,0.00358316441939155,-0.0111164239381675,-0.0161722132702661,-0.00919540943321462,-0.0320855705109503
"1098",0.00476044459550429,0.00324177980084173,0.0028760647983519,0.00292715873578753,-0.00632739503411139,-0.00220458864353357,-0.000162943837989649,0.00547924471999073,0.000341224255415495,0.00103589746505772
"1099",-0.00769918359203248,-0.0159244250784273,-0.0210324184661549,-0.0218889581873297,0.00902108219077524,0.00389364968316985,-0.00912503915975116,-0.0118899770380899,-0.00654881660546602,0.00172481566061466
"1100",-0.00634124797449243,-0.000468939868672247,-0.0058592836121425,-0.00149175833209736,0.00557391065760937,0.00241063011832221,0.00230213543822622,-0.00200546149119241,-0.00178541503174445,-0.0130854680616797
"1101",-0.0001498833508502,0.00187716257226622,0.000982250721778932,0.00320158208867682,0.010249630637972,0.00292878798071206,-0.00147624252733347,0.00728445674159506,-0.00433370036230651,0.00244246696417449
"1102",0.00893570210593087,0.00702544099644564,0.00785077780314869,0.0161702146563503,-0.0132513982686521,-0.00573574197425097,0.0111729372618266,0.00798003652198287,0.00594169524866328,0.02018793134022
"1103",0.0023815008964827,0.00837232414580158,-0.0146056315968759,-0.00649087764494194,-0.00042005369854814,0.00104899072705344,0.00194987776565858,0.00569052618336752,0.000343324161676151,-0.00784711418311368
"1104",-0.00794455737260547,-0.0161440442566538,-0.0108695913372827,-0.0080083036605606,0.000525048400613626,0.00240940278197943,-0.0102173232338905,-0.00787233903533813,0.0126331004174296,0.00928471077985238
"1105",-0.0116011288018688,-0.0241444914315502,-0.0149850855705557,-0.0208199700056262,0.00482559237083757,0.00135897340017954,-0.0104865119978585,-0.0176051144187829,0.00230522061478,-0.0160136901516122
"1106",-0.000832884022130886,0.0031229427331243,0.0121704024885467,0.00998043824937489,0.00375811089236011,0.00104368049909631,0.0029803276032927,0.00555327138047446,0.00514099972751136,0.0135042207483271
"1107",0.0033345313941533,0.00933903292775318,0.00200416067562226,0.00214823051318169,-0.00467977702144318,0.000104916361312934,0.0041274247856371,0.00301216819241645,-0.0000672589021404324,0.0181072403749749
"1108",0.00460773902644496,0.00972713817478632,0.00899975779770656,0.0128620132868975,0.00856907993775913,0.00552493255986741,0.0129894310814249,0.00725703166335623,-0.00242294383600838,0.00369129388523048
"1109",0.00383440395944112,0.00798887292519312,0,0.0105818673084028,-0.000414148248295887,-0.000104230124897464,0.00178544062297137,0.0111801931601296,0.00998513014448021,0.00568367458562014
"1110",0.0104113185094477,0.0219113620156455,0.0178396004296768,0.0163348840889042,0.00228028253755208,0.00155610376581516,0.0174984471516797,0.0122851745579813,-0.000400788251184836,0.00565158721344039
"1111",-0.0224610030094441,-0.0278284684496696,-0.0126581764643997,-0.0179271148431203,0.013514793546656,0.00824079472272188,-0.0281848771082275,-0.0177186389694249,0.00180436381852678,-0.0125619145801649
"1112",-0.00106154150502735,0.00821223626064316,0.000985982793067164,0.00944199528395639,-0.0190500290236005,-0.00597108343718156,-0.00573477605406225,0.00716573859243619,-0.00273500092762313,0.00870430105841091
"1113",-0.00994471803159769,0.00744684886581859,-0.00886695828912032,-0.00498859457119549,0.00574268798706834,0.00393521329524837,0.00362558644994149,0.00147197248277409,0.00481606020066883,0.00398275562528294
"1114",-0.010581207080948,-0.0157080400245176,-0.00994033862932375,-0.0160851863565665,-0.00757827001037892,-0.000618600982531192,-0.0142857741725494,-0.0100441518885171,0.00173076153820562,-0.0115702605873167
"1115",-0.000619725855958819,0.00938746258080858,0.00803230466745508,0.00785551789345917,0.00460303719486244,0.00185835004981949,0.0119941821238081,0.00296940387539357,-0.00039871080273024,0.00936459327804839
"1116",-0.00418732037627645,-0.0169729318630751,-0.000996034001490065,-0.00716244882786965,0.00780883514580299,0.00216353312658502,-0.00477382054968745,-0.00764856180035567,-0.00405531184756425,0.00828362085452339
"1117",0.0076311267808078,0.0130087226140259,0.00697907406370968,0.0078508019740835,-0.00402943559039937,-0.00400976086687388,-0.00926247582366124,0.00372969723987526,0.00500634143256584,0.00558665132076031
"1118",-0.0139105251059427,-0.0263832291115101,-0.00990096909755545,-0.0216841763456169,0.00767656978018083,0.00320028935389893,-0.023705927331904,-0.0173395217731898,-0.00876722248628092,-0.010457541356911
"1119",0.000783592270041877,0.00263774852166376,0,-0.00172166303867116,-0.00504442801248639,-0.00216073687789042,0.00188097783982721,0.00252082981845625,-0.00984991256198364,-0.00660506552415063
"1120",0.012686072416406,0.0141114533035773,0.019999986103622,0.0150894529840728,-0.0151055624198898,-0.00794011516166127,0.0157019525461761,0.0145838478820521,0.0060905053504634,0.00698149320234909
"1121",-0.0177852904303801,-0.0360847820494319,-0.0196078297804899,-0.0214480667383177,0.0181740768093566,0.0108094225125173,-0.0164674560667873,-0.0195786270177615,0.00302681782507319,-0.0267415394978376
"1122",0.00220458306840654,-0.000489601589313549,-0.00300017017273246,-0.00759578437576225,0.00453965375816234,0.00277658399419534,0.00700477801886046,0.000505446461664505,-0.00100586108522871,-0.00407053551353975
"1123",0.00298408852094156,0.0124848407259399,0.00300919827965496,0.00131216233341558,-0.00472479839567086,-0.000717650229067224,0.00848306679282529,0.00319167432753953,0.00651138479887625,-0.00442780233597684
"1124",0.00511593112879072,-0.00362674958240083,0.000999902320041102,-0.00152859810613448,0.00123829348242066,-0.00153896291474731,0.0105991162301788,-0.00254536102855052,0.000600220080029246,-0.00547389412708488
"1125",0.0137039361337852,0.023268356752534,0.0169831528955764,0.0183726136539146,-0.00443213712318857,-0.00133623157754903,0.00882298002968596,0.0130137971377968,0.00486566689905787,0.000688055927610343
"1126",-0.00602550800756818,-0.0126058245569975,-0.00118920050325444,-0.00995686419982011,0.00062117969618658,-0.000412052030239862,-0.0021450953007387,-0.00881619966269309,0.00152566998957515,0.00446882846379237
"1127",-0.00287553483815173,-0.0122758822777612,-0.00198418031403391,-0.00131447792026018,0.00765692169782062,0.00525050683214467,-0.0183561437857297,-0.0030497276034549,-0.0175508902062754,-0.021218265704642
"1128",-0.0116136355750723,-0.015660184952209,0.00596426122081617,-0.00175527806941889,-0.00421001164559009,0.00419970010644488,-0.00108806399188743,-0.00994126899727477,-0.0140218488343495,-0.0118882007975992
"1129",0.00891138589778073,0.0111112010930867,-0.00494051815345331,0.0116482996304228,-0.0137141993301614,-0.00387605280015824,0.00527589391578021,0.00437679139217018,-0.00362367713741552,-0.000353779382827213
"1130",0.0130528416882365,0.0119877730667293,0.0119162179561645,0.0136868139232353,-0.008050210712503,-0.00921445395676757,0.00829515197306652,0.0125610057668513,0.00349968444382576,0.0176990911858448
"1131",0.00856412213485935,0.0194968171969947,0.0157019522503108,0.00921544021879805,-0.0066402626973604,-0.00599354555417853,0.0110811682804304,0.00911427953361854,0.00642770765769596,0.0180869597716493
"1132",0.00956229492484617,0.0186395402749577,0.0077293705126138,0.0108304122607257,-0.00159149863529862,-0.00343070336133611,0.00132813565251655,0.0130455991429668,-0.00801734648811947,-0.0105910798016576
"1133",0.0147762291627347,0.00879270252605791,0.00862906297534383,0.0117647447970159,-0.00159937461467785,-0.00249895789974475,0.0179107638906659,0.0084198958532602,-0.00732881506849314,0.0013812676985363
"1134",-0.000821489588575974,-0.00777390673119005,0.00190108243814024,-0.000415273945415739,0.00224303386618496,0.00628974152016859,0.00619087456053657,-0.00736749162701977,0.0186297669937789,0.0134482335920072
"1135",0.00119597367187829,-0.0104461849659895,0.00569253446459528,-0.00664721841236771,0.00511476519428045,0.00177089777194439,0.00615287348030269,-0.00395862098680566,0.00867031739245672,-0.000340247139329009
"1136",0.0103751015384659,0.00791709086266801,0.00660382929499281,0.0138017262500372,-0.00296814899789477,-0.00384743683120414,0.0125521068520591,0.00596107867827111,0.00161164457426244,0.0211027479228436
"1137",-0.00709206748062241,-0.0147579933494356,-0.00843496937906552,-0.0113450251687184,0.0141426258334869,0.0106482252132893,-0.00349620246514404,-0.00691311345379286,0.00737516623701651,-0.000999986380040063
"1138",-0.0180804219042239,-0.0374487355632307,-0.0122871366012334,-0.0279573486178677,0.0149947802128694,0.00764375802295425,-0.0188199868322678,-0.0236202606488154,0.00891844259567387,-0.00767430506191968
"1139",-0.00431912459170702,-0.00803207575528686,0.00287046445194217,-0.0100881062132717,0.00340859966630092,0.00143521708898087,0.00341382351215946,-0.00127312718709127,0.0077842076069452,0.00874238413852768
"1140",0.00334854099356652,0.0156879929317106,0.0190841577183118,0.0162620135150546,0.00278000924182953,0.00163758357269495,-0.00842408423922114,0.010454097329742,0.00896769630247563,0.0136667549848453
"1141",-0.006902358882513,-0.00722474745085999,-0.00936333276783263,-0.0106677930545386,-0.014270940947953,-0.00572324421011627,-0.0111092118132753,-0.00782261687782315,0.00259500455816153,-0.00559029126745914
"1142",0.00580471313424114,0.00150576541052416,0.00756153184877251,0.00625409791194675,0.00166627780823658,0.00411187117598422,0.0109037540238022,0.00508635468183605,0.0042707650439715,0.00892861944212275
"1143",-0.00820096874225418,-0.0175393829032303,-0.012195220452093,-0.0115732324459762,-0.00967030072455621,-0.000614410881066396,-0.0089882341972759,-0.0129049678513561,0.00882738419125095,-0.00557203579296839
"1144",0.0162314346071102,0.013261803705414,0.0123457799603628,0.0145275735175312,0.0207891835356904,0.00379033227449077,0.0173153270375774,0.0115356100864843,-0.0121990350297424,0.00692156308141456
"1145",-0.000602816548436635,0.0135917863134498,0.0103189974824847,0.00299187694902336,-0.0118286448735961,-0.00489812835629677,0.00745658900683033,0.00608229230102464,0.00879348225026555,0.00327327776015629
"1146",0.0138714066777867,0.0273154752217561,0.00835654336295133,0.0159812322476318,-0.00770242165940949,-0.00553763488245218,0.00643593468100323,0.0118384021752265,-0.00762723990187819,-0.00489389755420977
"1147",0.000668947453526414,0.000483780140561718,0.00184166997740198,-0.000629081064465908,0.00755268645403961,0.00381536979715458,0.00511567152594794,-0.000995627492246465,0.00833167334067442,0.00819671052420667
"1148",-0.00557276039417098,-0.00579858747604145,-0.00367664806566648,-0.00209864361516776,-0.0109315753510808,-0.00318477407156459,-0.0112929598635145,-0.00647875828146005,0.00781450832098751,-0.00487801563658707
"1149",-0.00373635911678527,0.00680408020364176,0.00184514755977849,0.00336503809614208,0.00684179134678353,0.00422507362023405,0,0.00476537978036551,0.00273298595990812,0.00784313079179988
"1150",-0.0204754657701758,-0.0263091952403322,-0.0165746862359859,-0.0176065650105628,0.000104154562266423,-0.00164189711111429,-0.0268660122897112,-0.0154767912551769,-0.00367625014448247,-0.00680941221417808
"1151",-0.00290954861027803,-0.00421442229673985,-0.00187260205799467,0.000853483962409918,0.00376377149067197,0.00195305990778949,-0.00148814677238795,0,0.000827056418003069,-0.00326472866915961
"1152",-0.00683463674067575,-0.00199110833499383,0.00469032857365881,0.00426342204434738,0.0197871485630174,0.0121052937093644,0.000496995347253781,0.00025374469117212,0.00616568749580604,-0.00818865621833109
"1153",-0.00425243051676172,-0.016463039969866,-0.00933707856948529,-0.00084885528527745,0.0100929640057161,0.00363754402434768,-0.0132385593848241,-0.00481615360514009,-0.00360093515197779,0
"1154",-0.0255476897915827,-0.0304338363178178,-0.00848237299129073,-0.0308052918460577,0.0300267608478788,0.00921216956726978,-0.0293479596215976,-0.0191035820118592,0.0240933488201032,0
"1155",0.00541881880716533,0.00706272238779238,0.00190108243814024,-0.00350729378792081,0.00196920446745041,0.000802464151709703,-0.00621949844427883,0.0111657602100885,-0.000185729316846794,-0.014861261469488
"1156",-0.0468414469948283,-0.0727272212342204,-0.0607211391418988,-0.0571930829228079,0.035580524967701,0.0132300892844357,-0.0483308842813005,-0.060605795709276,-0.0052635207980829,-0.0378813261809202
"1157",-0.00149659123836232,0.0240895817848013,0.00909090724606343,-0.00653287660814927,-0.0288531273301255,-0.0115732608506508,-0.0206431899294298,-0.00328066614341971,0.00690986682588313,0.00418112739105347
"1158",-0.0651235560366372,-0.0820570123974501,-0.0480479330447384,-0.0833728603073269,0.0315673202266933,0.0159125108397875,-0.0850587205780318,-0.0811849810080102,0.0331993508500772,-0.0371269529125423
"1159",0.0464995743294172,0.0694277232257374,0.0515247177170461,0.0586729655249294,0.00303172962698972,0.0058118460666845,0.0925583365822567,0.0800002835662712,0.00891578533137238,0.00972978201500774
"1160",-0.0441779872230738,-0.0696571991621485,-0.0460001698497129,-0.0530009759174319,0.029753795487051,0.0132222749973778,-0.0235116316850145,-0.0527915801144304,0.0354071583215281,0.00428252295001075
"1161",0.0448836836344544,0.048817021620561,0.0377359035491276,0.0552010061426156,-0.0504497893492691,-0.0146928005334548,0.0466272791978992,0.0469795833059219,-0.0219383775697288,0.0216773984576242
"1162",0.0067332473089381,0.0251286647503308,-0.00909093623649715,-0.000484689039714103,0.0198032855635211,0.00696566561022594,-0.00146059896663941,0.00780401227288441,-0.00456807613469989,-0.00139135691917081
"1163",0.0211648648155069,0.0239551653465975,0.0122326283018299,0.0232614448168864,-0.0101351637042607,-0.00370237644752147,0.0356554248856416,0.0210175289176395,0.0107666175750627,0.0121908874330814
"1164",-0.00853924073719281,-0.0174100824313808,-0.00805661003568603,-0.00852474394546665,0.0165550079313546,0.00459585738250246,-0.00370748537729249,-0.00839638689102373,0.0123399008322485,0
"1165",0.000669061258789627,0.00664447485273034,0.00101538689349612,0.00716497595169008,0.0175090230592452,0.0070086563718621,0.00124039448062163,0.00655552384164948,0.00287488503765965,0.00860291493408494
"1166",-0.0431184500151818,-0.0539054639712606,-0.0344828670230404,-0.0471894790841524,0.0205385068147403,0.00522016782221235,-0.0430091111676215,-0.0331071735123707,0.0189198660580194,-0.0245650104809031
"1167",-0.0163309049859958,-0.0200579922385654,-0.00945365889541538,-0.012444433144035,0.00806792118760868,0.0010578797180365,-0.019974174608226,-0.0117876415105533,0.0125478054661952,0.0178383776501641
"1168",0.000799442077776158,0.0115690962027457,0.00212082580451778,-0.00100789270096968,-0.00251766612726612,-0.00182506071881394,0.0018872030680448,0.00369195881334106,0.025784935133953,0.00171818966189541
"1169",0.0329102755787292,0.0340177915627853,0.0190477353248888,0.0350656338505093,-0.0137939642034028,-0.00404189185737791,0.0246750300288998,0.0271649673367291,-0.0374884779779724,0.0102917024523768
"1170",0.0140844901476018,0.00425406610530299,-0.0114228086732449,-0.00974914593582077,-0.0284305474773445,-0.010725680979052,0.0112136334609632,-0.00110212122024966,-0.033883064489031,-0.0101868622966957
"1171",-0.0152437833084482,-0.0276760515469363,-0.0136553319674453,-0.0194437223257118,0.010820469946426,0.00615305544935074,-0.0210873577991962,-0.0170986924652575,0.00413636484018753,0.0044597718600301
"1172",0.0145336414845993,0.0116181493531595,0.021299090926902,0.0170684399258203,0.00986681953424928,0.00320382127900443,0.0148558899632005,0.0134678848350405,0.029647249769974,0.0112705134484055
"1173",0.0287363594391352,0.0267008501465476,0.0135558978137826,0.0323295275883317,-0.0138258797929125,-0.00657987970922802,0.0318393283597294,0.0271317829457365,-0.0201724346640422,0.00337722592734591
"1174",0.00263673051750657,-0.00782967652843281,-0.00411510045154917,0.00143443438424518,0.0160760151322974,0.00691561318126221,0.00390135986539408,0,0.0299615103223965,0.0134635385750419
"1175",0.0044379574956821,0.01944739178771,0.0175617256936811,0.0205300588284778,-0.0154536621392429,-0.00357908488999958,0.0107755915388013,0.0150945956730049,-0.00770522028904908,0.00166055506291896
"1176",-0.0104730111683566,-0.0102295294945577,-0.0091370542993352,-0.00537992280072097,0.0211979232990853,0.00796931856958882,-0.0167776939277996,-0.00929384611503958,0.000843990542178652,-0.00696293982860552
"1177",-0.0255498401220666,-0.0270947793953504,-0.0163934136987397,-0.0225777106262481,0.0324859444239283,0.00917041179076805,-0.0241735222112927,-0.014473257572681,0.0301906457016543,-0.0053421641792456
"1178",-0.00729752940036354,-0.0422051386666875,-0.0218748561236467,-0.0103467664955715,0.010399431797071,0.00133941780747748,-0.00218531887949347,-0.0190375569964789,-0.00185555004760019,-0.00335688875632811
"1179",0.0282076651043153,0.0305756100419607,0.0191689862182767,0.0296621486805764,-0.019088998750286,-0.00534981703007786,0.0335886298869545,0.0202383654977429,-0.0318206243352855,0.00909395082323083
"1180",-0.0103915629515221,-0.0206517231285799,-0.0125389249133422,-0.0221961307888237,0.00896778812728094,0.00489774953898592,-0.00724131596074162,-0.0187497087883136,0.0267110681419576,-0.00667547638088173
"1181",-0.0262097448481103,-0.0380158716128733,-0.0232803190551093,-0.0338079832378504,0.0106659491390646,0.00487412662227005,-0.0281087772592492,-0.0288010651189249,-0.00610528030477187,-0.0157930705888282
"1182",0.00647007204206984,-0.0101883223583247,0.00975080886193846,-0.0019995193006842,0.00105498362985057,-0.00304330672746367,0.00311191483817908,-0.00228114573839189,-0.0223021531096097,-0.0023899317720053
"1183",0.0091711932018923,0.00842159401424514,0.0171673481398888,0.00150268919148289,-0.0142313932316485,-0.00295691740372783,0.000912472938386921,-0.00342942877121999,0.0105846777674159,-0.00308004014999508
"1184",0.0138438094186717,0.0238169133263189,0.00421928000795857,-0.00275093183946484,0.0084662957764341,0.000573892786457808,0.00565188585043153,-0.00372809400269014,-0.0074492329570105,-0.00480608216168577
"1185",0.01725761417982,0.0259819762392925,0.0115547969075782,0.0145436678622164,-0.0152884331952591,-0.00745900154768631,0.0193978679146563,0.0146802415537273,-0.0158569656847878,0.00413940847517402
"1186",0.00591839183817511,-0.00294454585329473,0.0103840463948299,0.00172992017473672,0.0072691686928481,0.00192732292392339,0.00818065927879696,0.0000861015792028574,0.00934635926650329,-0.00446586426941942
"1187",-0.00995703424799366,-0.0318962465873753,-0.0143885221009118,-0.029607399260973,0.0190661626812123,0.00817319279911133,-0.0197565206235537,-0.0234690362128591,-0.0154519173746062,-0.0169082305750911
"1188",-0.00116374551964393,0.00671152259306584,-0.00104255648161067,-0.00737332514995159,0.00419678004852764,0.00133610310277654,-0.00287921891646914,-0.00175825253309592,0.014251924461969,-0.00175497785306811
"1189",-0.0294583174868408,-0.0300002110760997,-0.0125261911009741,-0.0371418599296489,0.0330841054952908,0.00428621147114416,-0.0478256314648122,-0.0258367031755106,-0.0124587723999247,-0.014767839573728
"1190",-0.0323243730988859,-0.0390501088542338,-0.0158562828078351,-0.0702311831279868,0.037585889141621,0.0092952414116505,-0.025208081439451,-0.0334537921007034,-0.0261535405531089,-0.0353319713791268
"1191",0.00602496688492793,0.0117033927232093,0.00322241272673307,0.0266096215917793,-0.0185997439471542,-0.00826974562454619,0.00803828316075594,0.00904236738750885,-0.054717538218559,-0.0177581084843996
"1192",0.0237802047710742,0.0285988908707724,0.0053533549517335,0.0150498241804933,-0.0160556630391001,-0.00416986666557517,0.012673130002651,0.0117431990235353,-0.0138923714538353,0.00338990068006195
"1193",0.0111835872971884,0.0296784177516356,0.0159742417827018,0.0318507792194807,-0.0153079201345693,-0.00666065866632004,0.0105888403151715,0.0186315690437824,0.0193552669202277,0.0168919313092548
"1194",-0.02041824673605,-0.018203920147383,0,-0.0300691488271239,-0.000341838764735813,0.000191717204101716,-0.0249570224408161,-0.0194903283076399,-0.0274544223540304,-0.0269472233298083
"1195",0.00790341150431439,0.0222496256105014,0.0178198107852805,0.013717404931886,0.00692124533557603,0,0.0148497360422215,0.0149849139766758,0.00947379330768272,0.0117601987558278
"1196",-0.0249892012759361,-0.0365779705657897,-0.0257466201507265,-0.0500678088725617,0.0251187631510412,0.00632102468664564,-0.026376650251734,-0.0343481067385027,0.00228282185699724,-0.0344957184688444
"1197",-0.0284576531742504,-0.0313773487719716,-0.0158562828078351,-0.0210825026107055,0.027520102593334,0.00926059209941199,-0.0470635947359261,-0.0190323009129241,0.0183475201612997,-0.00504847487959281
"1198",0.0219226292073293,0.0223517129764317,0.0128894659411198,0.0154250184219995,-0.0126805807977467,-0.00510293053511568,0.0377670967062185,0.0104958278319489,-0.0206262913495028,-0.001951653922452
"1199",0.0185153043031305,0.0186947333303038,-0.00424177335039622,0.023215793931284,-0.0071986757744017,-0.0041789202898973,-0.00759827328820151,0.00629541633057418,0.0115453438946038,0.0140790482234632
"1200",0.0180913027214769,0.0339034900469624,0.00425984263737234,0.0330532528238641,-0.0184576367830029,-0.00696258947698825,0.0276042546591879,0.0272129391653921,0.00645928731208456,0.0208252518572627
"1201",-0.00669578582098251,-0.00842364622700331,-0.00530226234100539,-0.0119308303515084,-0.00738770465335248,-0.0051863227168456,-0.0282352347305876,-0.00243601372569813,-0.00816257685330624,-0.00453344997004712
"1202",0.0334456500373508,0.0445992424107975,0.0255864277962827,0.0447310838894011,-0.0141237794598774,-0.0105233292939787,0.0482241729978263,0.0335773299902065,0.0256942529203403,0.0223909381486429
"1203",0.00100339130349969,0.000290647473973227,-0.00831623061510023,0.000525463694717621,-0.00334591472088663,0.0033171756684256,-0.0184791646928353,-0.00797393352080156,-0.00716603155102513,0.00742391804903431
"1204",0.00877206637931471,0.0223577090418623,0.0062893573707401,0.0280914850263596,-0.0145460004286414,-0.00340363507928709,0.0162776805324054,0.021435022224614,0.00715600837177011,0.00184234981324116
"1205",-0.00198747567328572,-0.00198807693040537,0,-0.00893793824138611,0.00995755239928275,0.0040012758024055,-0.00694716317447286,0.0046631499694898,-0.00588014228470357,0.00220658761071491
"1206",0.0170938939477643,0.0133750394800765,0.00208350897459586,0.0200979710084426,-0.0145296203280771,-0.00495681853989116,0.0231248832150841,0.016536369236966,0.00677751681865324,0.0227523610500662
"1207",-0.0190910924239078,-0.0292051276453844,-0.00415799597064914,-0.0338468518147245,0.0172880769365995,0.00654425563745042,-0.0229820237317261,-0.0231163897393127,-0.00477355586683803,-0.0143524120639776
"1208",0.0195458583589714,0.0161989840077379,0.00939444859357086,0.0266667835571976,-0.00621094394354171,-0.00106729088951951,0.033048061505681,0.00964061646328052,-0.00479645199841494,0.00546057776377684
"1209",-0.0118290356587801,-0.0170794534139643,-0.0155119378762678,-0.01909873897376,-0.000347005686427315,0.0015538997647877,-0.0124199981537663,-0.0144675711252096,-0.0121725225450452,-0.019551117232251
"1210",0.00437547202542121,-0.000868711191681637,-0.0031514507635183,-0.0192107843886713,-0.00712064978150284,-0.00203654693194255,0.00609765365121806,-0.00411056783397512,-0.013135616849178,-0.00147700870732781
"1211",0.0189874416773179,0.0315941239323667,0.0105375722057368,0.0285865461535773,-0.0105826369202024,-0.00184674159919207,0.0295458878563095,0.0250591972398599,0.0110920958080218,0.00517744365051964
"1212",0.0122606562624383,0.0126439003868388,0.0104274502523896,0.0391145959368775,0.00167963517983094,-0.000486775144937557,0.0264896204012282,0.0132296343593021,0.00940320939309913,0.0158204292876116
"1213",-0.0194435013062375,-0.0174804823164756,-0.0144476820988056,-0.0198117167938078,0.0254148035423789,0.0085725965812613,-0.0154124748669466,-0.0218562776634258,0.0283815171188295,0.0032597558763543
"1214",0.0101586233839941,0.0180740895736806,0.00209393631205934,0.018444105860016,-0.0174696786190189,-0.00734080311484642,0.00928320048124531,0.00783491176355144,0.0109305999379332,-0.00577620555844283
"1215",0.0348348732482655,0.0590845862379499,0.0386627997818878,0.0607784842139563,-0.0338974891103557,-0.0120658759946684,0.0427411548646173,0.0457819375357957,0.0128435428737232,0.0265069102104287
"1216",-0.000233233596525273,-0.012571910428561,0.00402413720052808,-0.00841888523715784,0.0105171023592316,0.0060079049952988,0.00311315077811525,-0.000826112713901095,0.000412810373114469,-0.0042447971617956
"1217",-0.0241056762811168,-0.0498676164839008,-0.058116294706786,-0.0375001994896522,0.0396554151560031,0.0134131677261893,-0.0131033494915647,-0.0338934797723023,-0.0134418056078823,-0.0152752847674487
"1218",-0.0278886107847377,-0.0424342981948428,-0.0127658119303212,-0.0242584179671652,0.0334743028325104,0.0119939296686993,-0.033717545351685,-0.0199658601260568,0.000239088089855066,-0.0119047844473724
"1219",0.0163116175916698,0.0134108408469942,0.00323261304913869,0.0306376339685102,-0.0124737031251556,-0.00239101068035064,0.0202494552231482,0.00407426764293572,0.0100369993417075,0.00620655986768326
"1220",0.0182272352828552,0.0322209605152979,0.00751886027025916,0.0102338861452271,-0.0137332936436103,-0.00469865066226127,0.0113411177186924,0.0133335856161327,0.0157340768453103,0.0123368135976034
"1221",-0.00609884463050081,-0.0167224088637601,-0.00213246749535301,-0.0065122850080469,0.00120293126273996,0.00298666327169927,-0.00753460405622552,-0.0051489156185226,-0.00506635799518773,0.00322572541378996
"1222",0.00621606592396873,0.00113410687438353,0.00854720929769748,0.00849721081592114,0.00635290798606336,0.0011522899251899,0.00247206225360475,0.00373803026996478,0.0241731920103063,0.0146481467086375
"1223",0.0128306944947001,0.0181198878908864,-0.00423728040599081,0.0117959673665695,-0.012796162455233,-0.00450882154412602,0.0119755365221628,0.0117444003510014,-0.00828664437733784,0.00492958259453546
"1224",-0.0369096871527755,-0.0631256576893618,-0.0180849663883224,-0.0585300297203237,0.020739949833968,0.00886647157867793,-0.0449004827711915,-0.0450171264356479,-0.0084134847485362,-0.0220743406300569
"1225",0.0094187056393884,0.0175125571083994,-0.00108356140610921,0.00657108030317,-0.0149002089226743,-0.00487182079847859,0.00091126476357295,0.00326128457171215,-0.00540482339842074,-0.0010748689279797
"1226",0.0188222771987185,0.030630036551083,0.0108461227080201,0.024102335974191,-0.00610177071242612,-0.00460808384123967,0.0258507742641663,0.0260048625308615,0.0164777843664707,0.00968441420898558
"1227",-0.00947420361251716,-0.0209452009080492,-0.00429183703497238,-0.013728782650488,0.0160830455786733,0.00626840088585867,-0.020053260302756,-0.0207373042787988,-0.00436887772716632,-0.0106571575633633
"1228",0.00494184178029711,-0.00578212799028122,0,0.00621426084491628,-0.00136149130348084,-0.0013414861569262,0.00869261035350499,0,0.000923810639557932,0.00718126704142441
"1229",-0.0158628155442115,-0.0180284912110713,-0.0183191921396191,-0.026926982225618,0.0091177327643277,0.00364683645346275,-0.00951527785877448,-0.0267646885072793,-0.0106714697123242,-0.00249550960909894
"1230",-0.0158770778446039,-0.0106604319183912,0.00109761416045773,-0.0253869753844794,0.00802269074484574,0.00200821205171109,-0.0179442368832305,-0.0163192057878079,-0.0257127230398438,-0.0232309291562415
"1231",-0.00106436812843991,0.00329250223066424,0.0043863667053925,0.00390684325443313,-0.000251345480781429,-0.00372197225274717,0.00719784327157869,0.00614446166612503,0.00311184309592405,-0.00146353550983858
"1232",-0.0190194910494835,-0.0256563490143351,-0.0196512723668243,-0.0321741255405037,0.00594933129399533,0.002778053118067,-0.0263881746099289,-0.0262594588995121,-0.0245793767026421,-0.00732866692535983
"1233",-0.00392786801374145,-0.00979793299897713,0.007795424597002,0.00348524849771525,0.0111617373241037,0.00305659483996212,-0.00282319361100447,0.00689856374930886,0.0110703241590215,0.00664450312592546
"1234",-0.0220656687235559,-0.0303029533759526,-0.0232043314777461,-0.0323267728544029,0.00980340969418414,0.00342786883157919,-0.0294449116942075,-0.0277172276194602,-0.00290361143189899,-0.0150348950280789
"1235",-0.00188759106212888,-0.00510213013964012,0,-0.0033133837661683,-0.0145212521372672,-0.00635856690896608,0.00350076315588388,-0.000640390919426581,-0.00867565359854827,-0.00819058292561925
"1236",0.0289667928999002,0.0503206608207667,0.0282808315503995,0.0479228342358173,-0.000496822691429366,0.0000960883110847632,0.0244180683007424,0.0326923325493607,0.0197675099057839,0.012387333873749
"1237",0.00284029337306935,0.00640808185321373,0.00440017807583382,-0.00449398142182245,-0.00819923881472007,-0.00191032371612054,-0.00283761431433471,0.00682795613564879,0.0015003300275962,0.0129774726077585
"1238",0.0411496956346142,0.0527594560236997,0.0328587718399855,0.0624004927082,-0.0156159985629325,-0.00583680862156366,0.0461013404561055,0.0554871307381717,0.0194750713244525,0.0117129078004778
"1239",-0.000159991910517188,-0.00576055245972518,-0.0137858090417977,-0.00299945919073985,-0.00501698714326682,-0.000289194885668809,-0.0101559473798399,-0.0175236016083975,-0.00293892896787962,-0.00361785859813823
"1240",-0.000880428933602739,-0.00144829636958244,0.00322590829218994,-0.00300815157916656,0.0140166672551771,0.00443717711528602,0.00164909108496314,-0.00356719374042003,0.00112009664799562,0.00871458986637008
"1241",0.0108923488104948,0.010443982091799,0.00750249522288549,0.0163440378365052,-0.00202344039893698,-0.000576440601902761,0.00932886900764052,0.0137233598174127,-0.0147214691847233,-0.00539956831462385
"1242",0.000316940903412277,-0.000574213811206703,-0.0117024268128887,-0.0136071743053483,-0.00954331615218107,-0.00259410936271742,-0.000725222712084306,-0.00706336967629473,0.00513976789398529,0.00542888193349578
"1243",0.00372240537047808,0.0066071975282127,0.0139936899598043,0.00401299075415307,0.0035815338472347,0.00452766508464153,0.00943059738905427,0.00533504905196991,0.00725413872505043,-0.00863930189363515
"1244",-0.0219363590003436,-0.0342466804055748,-0.0244162016032691,-0.0359729195391156,0.0124902796964859,0.00508326198201292,-0.0238950429676412,-0.0341979511289979,-0.0201888909157812,-0.0127087255023969
"1245",0.0169422314072345,0.0257094522084074,0.0228511536225338,0.0202123264768743,-0.0205605576278078,-0.00687050028754732,0.0198787337805584,0.0149575165317801,0.00253041336378867,0.00367777219365739
"1246",-0.0145974849583087,-0.0342842273410426,-0.0170214591409811,-0.0375919847856779,0.0111389688267027,0.00345871664385711,-0.0178668090293056,-0.0315792886523882,-0.0265023386959977,-0.0128252236904338
"1247",-0.0093388668576373,-0.0167064117643142,-0.00432887295767659,-0.00923723625875261,0.00932107312210606,0.00459606382136846,-0.00882039362077702,-0.0102483471520022,-0.021853249526105,0.00408313009436156
"1248",-0.0106461760764095,-0.0109225700369922,-0.0108693275156944,-0.0143847151799757,0.0188898011760008,0.00419341279690122,0.00574707617834069,-0.0128648659773571,-0.0350899217751327,-0.0354898435017028
"1249",0.0036143252152836,0.00429476628357617,-0.00219808161287094,0.00648648451990286,-0.00370752992579837,-0.000853837791060519,0.0136403730605337,0.00985375291697355,-0.00366274448075565,-0.00498276289883115
"1250",0.00148269635469278,-0.00763588869252729,-0.00330394320961391,0.00751883776014362,0.0116614797702008,0.00484462892638904,0.00836541681170688,-0.00331914809125033,0.0190375760646284,0.00808941651852191
"1251",-0.0106916676331393,-0.00447568431570322,-0.0143645680310085,-0.0258528322586505,0.0126715291764228,0.00340304249255952,-0.00973840810169435,-0.0150495374910073,-0.00231914584343618,-0.00458549768908145
"1252",0.0302601719559332,0.0384012889783405,0.0256408655886358,0.0419024577295903,-0.0249456355484006,-0.00904464753446288,0.030231120373363,0.0367361961029471,0.0136243369801878,0.0230327116103957
"1253",0.00193626271214309,-0.00541171286194719,-0.00995574353675388,0.0031813047673428,-0.0139096508986717,-0.00323271792836444,0.00141412560021936,-0.0119161868939609,0.00114669387556865,0.00712943567986613
"1254",0.00885909084964576,0.0120918737250855,0.0067039575247978,0.0132137257740863,0.00419861847398795,0.00124067055151889,0.0136810434167058,0.0111078263284374,-0.00712656510240339,0.00111779615846253
"1255",0.00894065021970314,0.00567498426534918,0.00776911021545001,0.00391227725239118,-0.0111206933689848,-0.00409678536982927,0.0049269703936099,0.00784672792470498,0.00173035767823948,0.00483808137586306
"1256",0.000791173834566949,-0.0026729634433541,-0.0121143357725916,-0.00961295067810497,0.00475028236540131,0.000565607280239799,0.00227641731607098,-0.00654004426350541,-0.00895652241003819,0.00444445986150788
"1257",-0.0131234929915058,-0.0157832368340466,-0.0122633668093072,-0.0167891918925264,0.0184887645198619,0.00632106697741808,-0.0108316969206752,-0.0163010392649364,-0.0250468329985969,-0.0117995140293872
"1258",0.0103339547043308,0.0160363422212768,0.020316074342025,0.0114730598211097,0.00182348652115372,0.00123741003987332,0.00830108478853409,0.0114723498327891,-0.00456864864310824,0.0029851108523391
"1259",-0.00491584109428689,0.00476470863053735,0.00774339094091769,0.00079110445869901,0.00322705817431723,0.00351725931206293,-0.00490481739671356,0.00283565447739131,0.0109751832107272,-0.00148807495388825
"1260",0.0159361319841949,0.0314166312569657,0.0197583959758065,0.0305748357038502,-0.0150104081735667,-0.00634712827341444,0.00616106183526011,0.0248189690415277,0.0258569173676915,0.0298061975373973
"1261",0.00156878492046397,-0.0103447860482367,-0.00107613371275805,-0.00562674497052351,-0.0118895529902459,-0.00314547608097615,-0.0111968884716953,-0.00367863857493433,0.00506675865914263,0.0075978046715317
"1262",0.00266244378208191,-0.0185829552812609,-0.0118537070789172,-0.00437259397330758,-0.00177986101813687,0.000191361989229533,0.00725444068984427,-0.0101538813487294,0.006827847311627,-0.0136445958527361
"1263",-0.0025773886204099,-0.0121304498027494,-0.0109049755661637,-0.0126580483847509,0.00789453080605163,0.00391991999666108,-0.00175667437410076,-0.00590585283240719,-0.00367601726249223,0.00436834231689986
"1264",0.00242767492677665,0.00509153742052315,0.00330786484082957,0.0104656418523008,-0.00176850615631108,0.000190321841627705,-0.00281521322508882,0.00250150409648509,-0.00445290720966107,0.00108748494039279
"1265",0.0086703104975161,0.0146008419225705,0.0120878002733418,0.0217502980458826,-0.00168742509110675,-0.00199991118443221,0.0111167278883106,0.0155957507263487,0.0136741150159743,0.0072410675824528
"1266",0.000542057347768132,-0.00616745899465754,-0.00434340153902912,0.000760482428306508,0.0130156505416128,0.00582030757224494,0.00890030675954079,-0.000614402437303929,0.00649268158404359,-0.00287566377870796
"1267",0.00239918435203879,0.0100472460926062,-0.00436188507683333,0.00405169871086031,-0.00141823620502723,-0.00208654381939732,-0.00657303066456139,0.0129072442943066,0.00444671515559247,-0.014059040274147
"1268",-0.00517315064258994,-0.0184317467224289,0.00219045064284362,-0.00907926433671713,0.00994213547998468,0.00446748218308457,0.00452737163520767,-0.00697814345848125,-0.00698347652501952,-0.00219379185917579
"1269",0.00388078225908317,0.0157972734793712,0,0.0190886778802386,0.00463294676235115,0.000946506362232702,0.00520017223500391,0.00824941354263742,0.00778604193727372,0.00696219963645928
"1270",0.0110561171380203,0.0184857551414892,0.0120219991407855,0.0252246956659283,-0.0121050120595538,-0.00311967938640245,0.0063803855258453,0.0139393686426112,0.00685361993769473,0.000363970964420313
"1271",0.00527636276963883,0.0164218706483028,0.00755948299156151,0.00876973465806841,-0.013753388827272,-0.00597582025107934,0.00633967777624767,0.0197248788081548,-0.00235151600180017,0.00436516390143638
"1272",0.00372734733315916,0.00255109104321161,0.0128617021266892,-0.000724584891686142,-0.0113256136258167,-0.00343396001801222,0.00476776247124255,0.0082064099363961,0.00527233590576648,-0.00724372798843753
"1273",-0.00257661755922023,0.00763351129595891,0.00423261305786959,0.00966657412428784,-0.00632588271275913,-0.0022022263461442,0.00305054520016723,0.00668608009709182,0.00672547018523906,0.0116745244053
"1274",-0.00113982514144562,-0.00280558117970198,-0.0094835990950668,0.00143599421100227,0.0018068793272219,0.0011509828333045,0.00557518604072693,-0.00779666923744571,-0.00704835113879987,0.00180315100471051
"1275",0.00836761866746216,0.00675253207889681,0.0127660461584185,0.0112335537851562,-0.00240432100033894,0.0047919933318914,0.012768578756444,0.0130967534450561,0.0272205612993197,0.00827933561250238
"1276",-0.00512979712434602,0.00251569031269283,-0.00210095404887267,-0.00401811466168123,0.0132561313105606,0.00534198187238188,0.00580658294188607,-0.00229853567551996,0.00510759530233873,0.00285608377297009
"1277",-0.000454833796802556,0.000557454502880139,0.00526327918843417,0.00522063198869671,0.00314340952615022,0.00303621402991539,0.00247384840299558,0.00518314095971451,0.0101631910046465,0.00356001051713029
"1278",-0.0034138308237992,-0.0153247317994962,-0.00628288436285618,-0.014400241155349,0.011772113536856,0.00340473118870266,-0.00871985177640278,-0.0077342671436087,-0.00556312951670035,-0.0102873049938557
"1279",-0.000380519062569418,0.00679143206520849,0.00632260858144496,0.00862289683904205,0.0115508120739762,0.00377105051569671,0.00514511133103634,0.00346443410482555,0.00761768141175789,-0.00250900001479271
"1280",0.00875713025889868,0.0207978573737269,0.00628276557974194,0.0220846936939343,-0.0114547503117944,-0.0034716351338252,0.00743061926718891,0.0161101318571222,0.00147658143614171,0.00323395006293814
"1281",0.00158537599774977,0.00220306595823283,0.00312187273055997,0.00278835344089257,-0.000419673605483561,0.00141605783565657,0.00213087749978458,-0.00141510227646768,0.00878747946198954,0.00250709217230694
"1282",0.0140183613623799,0.0189558661749092,0.0031119216243265,0.0166818631322894,-0.0214885907301468,-0.00791909399427471,0.0143931686229317,0.014459500143422,-0.019935714353656,0.0117899484229973
"1283",-0.000668757610198911,-0.00620100680608915,-0.00310226761066446,-0.00843192820911376,0.00995055483072593,0.0027554200171469,-0.00483713826027177,-0.00614882195952238,-0.00274401099226917,0.00494350813762146
"1284",0.00252876860170193,0.00678231922439765,0.0103730916934424,0.00206840104522166,-0.0124011316684053,-0.00644388687078867,-0.000810126691695334,0.00337458576597416,0.0150735979514007,-0.000702731107745658
"1285",0.0029676145439379,0.00323361627290297,0.00410682448898214,0.00711024471247157,0.000773994235103714,0.000476740508100315,0.000648644478252747,0.0053253445357635,-0.00707128474492547,0.00457096435919468
"1286",0.00125756375389408,0.00268610279935566,-0.00306728861869998,-0.000455779826920688,-0.00747677271168856,-0.00228809528439222,-0.00729223341975005,0.00139366282730924,-0.00284864094955495,0.00525029928143272
"1287",-0.00738758479537305,-0.0192876606530892,-0.0123076304650366,-0.0221003337761296,0.0129880323853702,0.00563775838483416,-0.0083251460181365,-0.0153114545703035,-0.00523750136323065,-0.00940102202020787
"1288",0.00744256739308469,0.0101065541264962,0.010383981561106,0.0163090728263446,0.00128228349616966,-0.000665231015402723,0.0113579607793306,0.00706813213816915,0.00221368913613551,0.00246042320711748
"1289",-0.00125598427359619,-0.0089235089235089,-0.0030830505522883,-0.00825301449791938,0.00529291807555188,0.00209190822200545,-0.00992815007651415,-0.00561508011853917,-0.00232821928028837,-0.000350626340403282
"1290",-0.00465989446758375,-0.00300159691194601,0.0164948594667127,0.00277392537120047,-0.00178328218964796,0.000759061557969343,-0.00493185450262923,0.00846987506230801,0.00592392310686707,0.00350749322354549
"1291",0.0110731125199781,0.0139573809003248,0.0101418453607813,0.0108344572487018,-0.00799673182121474,-0.00455095925062521,0.00826028721990379,0.00895852762020599,-0.000654339416725214,0.00454391175146429
"1292",0.00264609433935648,0.0043182878640744,0.00100397078131831,0.00182431109830894,-0.000256917873996731,-0.00104741323297519,0.00163857183561333,0.00721422898096846,-0.00386901190476185,-0.00173971176077381
"1293",0.000439988815700065,0.00134370530903904,-0.00100296383493326,-0.0040972524571673,-0.0110658955329556,-0.00362351946066619,-0.012432622564333,-0.00688713438172572,0.0219300739074966,0.01568487205973
"1294",-0.00322447091431599,-0.0050990578489738,0.0030119692906807,0.00182867127329756,0.0125772885044135,0.00392315988264835,-0.00811643761730896,-0.00693472421921504,0.0112267451473103,0.00926559358588586
"1295",0.00441083532587916,0.00971114525856986,0.00600604786318049,-0.00182533333865698,0,0.00142994754916725,0.0116900565833686,0.00810044240784658,0.000462599740226777,0.00306014184494452
"1296",0.00219550375245858,0.00854923570499344,0.00199024225393507,0.0100569981186751,0.00651063025454923,0.000761601633840092,0.00280607035350178,0.0119148593470249,-0.00456599226526433,0.00610175144674652
"1297",0.00167991048268679,-0.00741721216950575,-0.00595844473763918,-0.00995686197650947,0.00885068106973375,0.0033289183649956,-0.00115243027002687,-0.00492883727903903,-0.00307727464616558,-0.00808621224280259
"1298",0.00291659464606209,0.00854061817055407,0.0159840316637869,0.0139430232148705,-0.00329004897044582,0.000474224090843078,-0.00758062037746643,0.00963121264491651,0.0104252069381223,-0.000339669258072273
"1299",-0.00392579021438655,-0.0108496052873783,-0.0176992088182166,-0.000676184218065257,-0.00609442944906624,-0.00397947453752923,-0.00132845782388791,-0.00572365297376864,-0.0530290606654832,-0.0037377712839286
"1300",0.00518136750008535,0.0136436623839418,0.00600604786318049,0.00947413930597052,-0.00941391968945737,-0.00323996695377582,0.00532105829793927,0.00986831471187855,0.0141214200429116,0.0156890517662007
"1301",-0.00304932548070025,-0.0113487751281974,-0.00995025184479759,-0.00245831123725471,0.00939180136161522,0.00401483081405196,-0.000330857961425512,-0.00488577330868867,-0.00162058098781237,-0.0100739096678047
"1302",-0.00407818302165508,-0.004003941409497,-0.00602985052335769,-0.0172487991709466,-0.00793853687272483,-0.00199943819789672,0.0081072167052596,-0.0043644105040016,-0.00414814245877471,-0.00474902210510297
"1303",-0.0146252455898338,-0.0399359964503607,-0.0080893000179334,-0.033508259345744,0.0121323405901037,0.00419788878199179,-0.0134579251456479,-0.0263015492964673,-0.0178086151937923,-0.0163598703524483
"1304",0.0069760126631877,0.0142380734803238,0.0061163372005324,0.0120283662996061,-0.00612134823860655,-0.00189981801563499,0.00432515576825665,0.012380167502583,0.00571609107036442,0.00450444281824036
"1305",0.00994887357234853,0.0253231536325937,0.0172238511915803,0.0209742298317772,-0.0100070242463897,-0.00295125544175523,-0.0023189403090027,0.0216789133194892,0.0100836885019957,0.00827878144789507
"1306",0.00386762660586282,-0.00697955952038265,0.00398413824371335,-0.000456521280128186,0.00198636335226388,-0.000763388941591558,0.00464902212631912,-0.00516880286239774,0.00665540904317163,0.00273687664164446
"1307",0.0000729090198803295,0.00162189852859096,-0.00992072122176646,-0.0109615692604759,-0.000172157783521421,-0.000287240685151846,0.00694083575944915,0.000547116308132978,-0.00787353023579973,-0.00136470329624794
"1308",0.0180257776313661,0.0178135031628575,0.00901819771477808,0.0272457132050588,-0.0175935953580817,-0.00716676548362394,0.0178893389152024,0.0177645355842053,-0.0167807831982463,0.00444138199630006
"1309",-0.00107112533967957,-0.00689435375724667,-0.0109236886218586,-0.0157339729339958,-0.0251955628625273,-0.0114543019264693,-0.00241864593483909,-0.00939861568321887,-0.0168206774463214,-0.00680273323384251
"1310",0.00578952485397766,0.00961281027826755,0.00803213640426526,0.00799263534092987,0.00153161416789227,-0.000292489177434518,-0.000646393741051909,0.00921639285596676,0.00946289987942417,0.000684922163946666
"1311",0.00138473875406198,0.00872768686346315,0.00597624973529531,-0.0011325548789618,0.00197775562832936,-0.000292222417004329,0.00598412657499003,0.00637937681385581,0.00136578716953339,0.0123204071609913
"1312",0.00392005431165132,0.00471948539726963,0.00297021874301184,-0.00385597609196009,-0.0119357347124049,-0.00613761188056561,0.00594844229682989,-0.00134308117402515,0.00179784869563826,-0.00169030813224702
"1313",-0.00291110662411331,-0.0117431751769635,-0.00987178217331175,-0.0173040634105102,0.00399642013914558,0.000489871827891397,-0.00239729885275108,-0.00995134001501607,-0.00903515710217606,-0.0121910687751201
"1314",-0.00163716164417549,-0.00580942994098665,-0.00498501811302132,0.00185344840426627,0.0113080945146191,0.00509474962894862,-0.00224295602115554,-0.00353143631727282,0.000499606554061893,-0.00239976354492633
"1315",-0.00720398032831349,-0.011420950456558,0.00100193040466778,-0.0152637138837692,0.00322018143176739,0.00126764354830344,-0.0118816049191763,-0.0109052951698383,-0.00399475670705129,-0.00790370781297056
"1316",0.00323303312008028,0.00698532089438597,0,0.00751531264627725,0.00945144790514196,0.00369972773607663,0.00406234833009789,0.00303172560134435,0.0122829599173986,0.00969855199605174
"1317",0.0140351423653315,0.0170758310782111,0.00700708895954683,0.0174826083987241,-0.00512327227670895,-0.00116404814600124,0.010333619221953,0.0129156704223692,0.0177675665063304,0.0044597718600301
"1318",-0.00310710885423726,-0.0115422959647333,0.00795229407247633,-0.00526921146169612,0.00719195076275247,0.0055356299857594,-0.000485085236763938,-0.00189902131374697,-0.00705589441809829,-0.00409837491775156
"1319",-0.00495872283813614,-0.0111467704919681,0.0019723535448064,-0.0168126403611232,-0.00141022432437587,-0.0017384327827461,-0.0022628885449798,-0.00679505140314962,-0.0105979536082469,-0.00960224010502808
"1320",-0.00170879891624598,-0.00778303269008052,-0.000984179686273512,-0.00117102311228512,0.00750317166426084,0.00416028474095187,0.000972099489840117,-0.00191573557992208,-0.00142403570751148,-0.0138504051469359
"1321",0.00413642521244606,0.0102786603360474,0.00295589479626401,0.00727001674528394,-0.0169104499862917,-0.00491392532897716,0.00841715358204653,0.00959693683344853,0.00520830856403953,0.0112359826673936
"1322",0.00731487608335302,0.0152609565133073,0.000981827964540827,0.0137369569146719,0.00554027150405401,0.00239552524953845,0.00642045136579394,0.010320449370306,0.00505802507580877,0.0128472255229006
"1323",-0.00408934744313461,-0.020833130241711,-0.0127573945941051,-0.00574198543754867,-0.0173288834496912,-0.00735385980591963,-0.00462526576196187,-0.01290322954037,-0.0187185648862335,-0.00445657267375199
"1324",-0.00991093801465026,-0.0258552689559963,-0.0228628066966687,-0.0180178963725313,0.013745984586131,0.00506910126388771,-0.0100945639377368,-0.0152503816123809,-0.0167614736178715,-0.0154959387610798
"1325",-0.000500211253981919,-0.0091236253856225,0,0.00541040526272418,0.00722582665691163,0.00446128237606369,-0.0043703959904392,-0.00359551064497488,0.00699695280848123,0.0038475546290011
"1326",-0.0112310422959893,-0.00446418523737035,-0.0061036905276256,-0.0147400475654865,0.0233811084932707,0.0102345686631542,-0.00959216990933842,-0.0049957432997626,0.00669570471474579,-0.00452973397957102
"1327",-0.0167850692159521,-0.0252243080852308,-0.0122826970358146,-0.0194728013399279,0.0113368569890471,0.00468340776316256,-0.0193693884842596,-0.0108786065966907,0.0108553118797552,-0.0133005924675427
"1328",0.00809408547148083,0.0169639268328183,0.0134715136150008,0.0108983693632969,-0.0119801996060828,-0.00390048221721917,0.0118846680723992,0.0118442816686399,-0.000186213525032453,0.0024831161464689
"1329",0.0130658536530768,0.0197907790473342,0.00511259232487116,0.0256346799699372,-0.00415653672553806,-0.00200532644394247,0.0142266783911766,0.0139357207273678,0.0101197611545394,0.0130927143080344
"1330",-0.0118883741870864,-0.0263376411996569,-0.0111901618088022,-0.0151833547890955,0.0161765990338454,0.00602858035929676,-0.00521923142105662,-0.00769668475313112,-0.011370565667558,-0.0101291689588564
"1331",-0.000656351778232533,0.0105350435304219,0.00205737429440145,-0.00498082074390671,-0.00145535184615608,-0.000285659952387163,0.0116413329017124,0.00332378082880846,-0.00242461290302975,-0.00988007454080853
"1332",0.0148123885094464,0.0208511069798401,0.00616029496647896,0.0114421358154058,-0.000600114268895613,-0.00104638166593374,0.00858971268614561,0.0124241609042202,-0.00130878094751663,0.00463293958054045
"1333",-0.0033799420130467,-0.00800426385435349,-0.00204089794416418,-0.00471366476542112,0.00291645414181341,0.00200014477352495,-0.00530283937443499,0.00245438101454409,-0.00586584711388449,-0.00957784323772171
"1334",-0.00642050133383498,-0.00528693460894625,-0.0061347802193088,-0.00449910321548197,0.00094083800839817,0.00114086087203424,-0.000484679994698034,-0.0043528096828428,0.000753217007761098,0.000358161290763714
"1335",0.00166994762989203,0.0125875148132877,0.00205737429440145,0.00689823205459028,0.000171009368322039,0.0000945135979075751,0.0105059469803126,0.00928990676437191,0.000689958005580582,0.00393840047884164
"1336",-0.00840873679832121,-0.0223755753006758,-0.0112933305971585,-0.0191355533462609,0.00726005916138983,0.00199402080204192,-0.00927725215751007,-0.0143474235897231,-0.00294588203974666,-0.00178321596697351
"1337",0.00380116381135709,0.00734667204270645,0.00623033592831779,0.0021677378288214,-0.00703894071073607,-0.00255797206314823,0.0127545862501697,0.0120842772195062,0.00144587910906413,0
"1338",0.0136919723349485,0.0165496541470023,0.00515984322393015,0.00913248214632767,-0.00512374019791617,-0.00123557882285441,0.0109994096082582,0.0108550722593397,0.00200873819192582,0.00571639657127987
"1339",0.00696894519271019,0.0066227008726909,0.00513355972773066,0.00619186979810071,0.0060085583335272,0.00332865377698499,0.00425746580846642,0.00375856551530052,0.00883350485006607,0.00213140957556313
"1340",0.00164094296728101,0.00520818715348192,-0.00306435818446671,0.00142024517741746,0.000853868814593817,0.00104344115297228,0.00486717628612876,0.00401158805418311,0.00217354531561553,0.00319035098056442
"1341",-0.00370400897509804,-0.00627189261221206,-0.00204926237770342,-0.00212717758902492,0.000255549578240588,0.000852150752360448,-0.00140632933370921,-0.00372940736309491,0.00309827726179579,0.00388694552119162
"1342",0.006219933299761,0.00768371518461985,-0.0102665953584101,0.00663142931494987,-0.00518649641524593,-0.00181956206954026,0.00876254258834797,0.00267374610764848,-0.00345934014518967,0
"1343",-0.00298421261402626,-0.0106207592448013,-0.00518692828762368,-0.00188214830567857,0.00704279740930946,0.00189885934388734,-0.00155136375836529,-0.00239997513208623,-0.00452523536029847,-0.0130235865097412
"1344",-0.00762548739349234,-0.0090834423099786,-0.00834194245807418,-0.00754346341545686,-0.000255740960468875,-0.0000947597191973681,-0.00341757806029219,-0.00908843029356721,-0.0100877703490323,-0.0110556673761554
"1345",-0.0161580602925778,-0.0172224263141999,-0.00736063863969971,-0.017577174661878,0.00784852174880823,0.00398035151009046,-0.00763842062201725,-0.012948561981894,0.00314524751119549,-0.017670375073744
"1346",0.000730250083980311,0.00819674544411231,0.0042372467644598,0.00362681492579564,0.000169261377125807,-0.000283102097241361,0.00565517083809408,0.00819889062781542,-0.00244559476738193,-0.00220261312828607
"1347",-0.00401194482551492,-0.0134567390961072,-0.00843894592525607,-0.0158998535536409,0.0053318313181161,0.0022662378267837,-0.000937428502108983,-0.0103008257318794,-0.0193613399627692,-0.00367920130409782
"1348",-0.00593163225705962,-0.0147769629821647,-0.00851040579899298,-0.012974483048442,0.000673495444242445,0.00084788884060627,-0.0023451584905323,-0.0106820347990967,-0.00980768589743597,-0.00775473278825167
"1349",0.00206282072677433,0.00519187970960644,0.00429143816809052,0.00421640099469545,-0.0029449702651021,-0.00141253110657269,-0.000940112004446436,-0.000276785842393545,0.00194214409307869,0.000372080552337062
"1350",-0.00301460743401671,-0.00487794120648877,-0.010683523668543,-0.0128426287987381,0.00826906960282314,0.00329929271239138,0.00423527858038408,-0.00498480216236363,-0.00781809115931786,-0.0074404513480204
"1351",-0.0110610100377431,-0.0204728873617209,-0.0107989857845252,-0.0227669734861317,0.0139747380315047,0.00441580544572373,-0.0121837464397527,-0.0125240948395484,-0.0145219850810365,-0.0131184545155544
"1352",-0.00574155686180877,-0.0156019594506337,-0.0131007105903591,-0.00870473395400018,0.00404418179767041,0.000280446461977446,-0.00490195973846941,-0.00930116154642602,-0.0105068193946103,0.00189894864774565
"1353",-0.0038246911501687,-0.00687807899270176,-0.0110617943502787,-0.0142046259009562,0.00287673944764411,0.000747778066700011,-0.0122356282133818,-0.0082501769063823,-0.0018698944213339,-0.0011372096858524
"1354",-0.0148310741621556,-0.0165613401065168,0.0089486811943067,-0.0136232144509609,0.0177035167222388,0.00373793320307536,-0.0276706711753603,-0.011761745003452,0.0223470884756483,-0.00227693068930646
"1355",-0.008558719627626,-0.00275562422834985,-0.0144125503521981,-0.00956175397065728,0.000241636428412795,-0.000651679824415385,-0.0102582161799133,-0.00725660159061448,0.0114528793562916,-0.000760813374248825
"1356",0.0171881630122874,0.0239484975494237,0.010123309457468,0.023867068097517,-0.00209332147025798,-0.00260846248893665,0.0205616274347382,0.0236840062855419,0.000646981546807091,0.0133231960579028
"1357",0.00174277946275336,-0.00329837850990267,-0.00111309381846691,-0.0104764505845661,-0.0111346860582486,-0.00214762684941139,0.00212958871902091,-0.00628401995600225,-0.0166181189764546,-0.0142750178179645
"1358",0.000529870159235335,-0.0105293280307589,-0.00780375375636477,-0.00688229851231248,0.00693558383571014,0.00262008576751982,0.00424946480865662,-0.00546112647773545,-0.003024769818191,-0.0110518353072266
"1359",0.00196539585015199,-0.00638513371548355,-0.00449468849517021,-0.0050636677956738,-0.00380844429589378,-0.00214629900985974,0.00309268880425839,-0.000867146683395048,-0.00138498223799577,0.000385351197087491
"1360",-0.00324435959206593,-0.00152988765638218,-0.00564321528067357,-0.0048219061492506,0.00374160286210001,0.0028997937970594,-0.00292073253790015,0,0.00838774827586697,0.00346682482868865
"1361",0.0121118333048746,0.00950047561552636,0.012485860502307,0.0282635278036116,-0.00307909223778635,-0.000839670999732034,0.0136698506087607,0.0138849649550634,-0.0108723413420644,-0.00422251234308701
"1362",-0.0145100872781933,-0.0258045756486026,-0.0134529437399317,-0.0172774115122138,0.0253615155295368,0.00952303432594293,-0.0232783107635557,-0.0199713097248801,0.00589325901487858,-0.0185043039401039
"1363",-0.0022009321456482,0.00124663432088945,0.0102273272562641,0.00426219469363875,0.0115745152706586,0.00388418926065359,0.00624568826606064,0.00378429669982094,-0.00190908427597691,-0.00864096828130689
"1364",-0.025177014213689,-0.0211641431203992,-0.0269967785366355,-0.0267903376331318,0.0237399294210376,0.00859020021482171,-0.0253183678059838,-0.017981500682194,0.0387811976909775,-0.0206023441985491
"1365",-0.000468019917911233,0.00699524913418226,0.0115607965464521,0.00436080666081362,-0.00790081302293311,-0.00576323392007749,-0.0070386348544601,0.00383969772928627,-0.00114281269841265,0.00566352009082416
"1366",0.00757234143554397,0.0031574357857429,0.0125712831486959,0.00271360172024693,-0.0133768055778205,-0.00331268396082951,0.019746785667538,0.00617819197272551,-0.00114421556058042,-0.00362030687199211
"1367",0.0224682327735801,0.0336794815837116,0.0158013484769939,0.029228656216727,-0.0199845817244134,-0.00655478623944505,0.0213505878783133,0.0362570683341776,0.00044551355762712,0.0185708895967318
"1368",0.000606268938169396,0.00182716848995401,-0.00666646163817064,0.00604791734863563,0.00151949257173833,0.00241644718143719,-0.00486143817821227,-0.00423253441678806,-0.0172381329389546,-0.00673799981177947
"1369",0.00795145633098127,0,-0.00894874463830775,-0.00862525052444796,-0.000239224580939057,0.000741390344912496,0.0125386332672226,-0.00510049915996136,0.00148864724919084,0.0031922947283809
"1370",-0.0126973949054925,-0.0112462681363305,-0.0045143737722364,-0.0145002577141462,0.0045519088887287,0.00268657357348068,-0.0196205204184768,-0.0150951510091079,0.00407164102815605,-0.0182974890606896
"1371",0.0114912141042007,0.0190595215836558,0.0113377413974922,0.0208666605454313,-0.00914271321733662,-0.00535833206695002,0.00935043408951231,0.0118561371045796,0.00708036813156299,0.00486217012124057
"1372",-0.00639496433730247,-0.00904987050920769,-0.00560538262726251,-0.00366879961400224,0.0098690304325344,0.00529444907118792,-0.00471347945351341,-0.00600184400303883,0.00421825367807882,-0.00766118603546284
"1373",0.0106003148773279,0.00700165174665401,0.00789179765816006,0.0071015651348687,-0.00127158965361096,-0.00267969754124808,0.0135533405311894,0.01121368496695,0.00400970608483031,0.0117837915331112
"1374",0.0102272496981684,0.0157193129592765,0.0145413333384934,0.0182814066227075,0.00556932888652018,0.00463214323751804,0.00628354065840941,0.0120371359062195,0.000570497622820909,-0.00160644505840102
"1375",0.00193831689140511,-0.00922620706164989,0.00220537871899129,0.00205195096251232,0.00537949687202377,-0.000276792974735596,0.0078449222293937,0.000855648724658042,0.000570178676385646,0.000804494238004771
"1376",0.009672670184248,0.023130189836249,0.00550030036382165,0.0161247594875984,-0.0130625157545399,-0.00341279713233011,0.00466373927761765,0.0170986896679863,-0.00487550835261552,0.00844052334810597
"1377",-0.00162126543708785,0.00703774436524318,0.00875277447287925,-0.00327435229046324,0.00494347670720652,-0.00203642729345244,-0.0012763288152936,0.00196134240010482,-0.00757192014324448,-0.0163411536663084
"1378",-0.0224386806273359,-0.0275945539306232,-0.0144548389171494,-0.0366220805818028,0.00531562680863917,0.00213369000918617,-0.0156523067244775,-0.0209730837503863,-0.0253253636896495,-0.0214749183216139
"1379",0.00770118862787639,0.0111042254999525,0.00666700061124326,0.00318541991386323,-0.0133374064639695,-0.00435011765640503,0.00081118149235393,0.00942575244783006,0.00407837773770869,0.00993788052228783
"1380",-0.0160342330886515,-0.0265405595701065,-0.0154527701620444,-0.0185234906933806,0.014557735451469,0.00548408860445448,-0.0055124956543835,-0.0116016181673529,0.00733750004807066,0.0102500893865118
"1381",0.00502555799894489,0.00626753714331851,0.0112108294768711,0.00862767929779129,-0.00394188869003642,-0.00221884058107924,0.00440189738001107,0.00973403873554068,-0.00741415216617314,0.00689934024072114
"1382",0.00901679277614997,0.0084087746584518,0.00776069645006561,0.00641543296342362,0.00158265687377512,0.00138962253927777,0.00633020358301328,0.0110572039325116,0.00137601236325557,0.00564301657149979
"1383",-0.00285357584814594,-0.00154421688393624,0.014301302392695,-0.00478080942116232,0.00244993390026238,0.00323836491854812,0.00838708541787181,0.00168288681206685,-0.0116469212635357,-0.0108217008893704
"1384",0.0249267398736965,0.0423755687483474,0.0206073625167946,0.0443020698938861,-0.0130073250463445,-0.00461112657619289,0.0227126430113198,0.029675056899255,0.0274081358343303,0.0433548923793641
"1385",0.00301244721245375,0.00919873054601927,-0.00318821209263942,0,0.0103177547642208,0.00463938413936282,0.0106351178286217,0.0103318419839615,-0.000644410069663981,-0.00194172110753565
"1386",0.00659274386890574,0.00793886465006532,0.0127931580728333,0.0199336954493066,-0.00768514628462913,-0.00249319229903833,0.00557111198672522,0.00430596232557101,0.0152815208016381,0.0280155820911756
"1387",-0.00451213472656298,-0.0239205878540124,-0.0126315605223641,-0.0105238531041365,0.0051100415849854,0.00268486974650362,-0.00461705401932411,-0.00911065953131807,-0.0113045466840351,0.00378503751243242
"1388",-0.00950321689858502,-0.0128510228128618,-0.00426407658837935,-0.0182323870145652,0.00929366050755509,0.00350928333143252,0.00139125360669712,-0.00432667584393021,-0.0126540730252988,-0.023001542465737
"1389",-0.00125497704664213,-0.000605568531430678,-0.00535371043379596,-0.00361130209659422,0.00881469333380602,0.00276030254344817,0.0020073632779305,-0.000814995556196574,0.00214680882813312,0.0177537984865639
"1390",-0.00872015403519599,-0.0042413238337734,-0.0107642979607504,-0.0111310505309794,0.00202843332830871,0.000458748572455869,-0.0118643610588545,-0.010328705342855,-0.0122695344448635,-0.0128934580304473
"1391",0.0001491287830786,0.00365098559631694,0.00217659142597859,0.00523550809382511,0.00124554401009069,-0.000916757365511334,0.00155928481448298,0.0107111697319091,0.00552094007969539,0.0111409573662571
"1392",-0.00484492156719429,-0.010306436106676,-0.0152010057799163,-0.0166664547702504,0.00707608444736429,0.00229515681023718,0.00435927520683199,-0.00624989889342797,-0.00261460871251018,0.00227960414753747
"1393",0.0167776998287412,0.0159267098827598,0.00992302401152001,0.0193325300154563,-0.00262505087210252,-0.000824187670800836,0.0108512591970322,0.0150394916046168,0.0101579595034524,0.0121305097542026
"1394",-0.00235726232006028,0.000602938215416904,-0.00436719305748223,-0.00233838962562882,0.00464528105183004,0.00219990537074444,0.00383334222423426,0,0.000454184510537026,0.012359496595415
"1395",0.00686691238164427,0.0042180242998735,-0.00438597950133768,0.0132811874123728,-0.0078603105345435,-0.00256091717548368,0.00840214954788276,0.00942937134953437,-0.00479868988009313,0.00110978658825989
"1396",0.00740713175442931,0.00690085679541297,0.00330405313311677,-0.0025699876669133,0.000543767423500263,0.00100851755554388,-0.00772619533835273,0.00400299369497548,-0.00273667816031353,0.00886924934503464
"1397",0.00262090305465112,0.00953508736428077,0.00768402762864495,0.00927616408397958,-0.00256190329002537,-0.00146590768456101,-0.0083966919536228,0.00318969132480551,0.00215617114362288,0.0120879356194799
"1398",-0.00914871902045666,-0.0242030009194759,-0.0239651238801355,-0.0148073616400825,0.0122189575039944,0.00394541915374891,-0.00338718737426846,-0.0116586426683781,0.00189068320867491,0
"1399",-0.0101118216710744,-0.022988519914049,-0.0133929609867391,-0.0261725927976761,0.00561265600333205,0.00164492699272123,-0.00602502441795671,-0.0131367047795918,-0.00416476220686868,-0.0209916867428366
"1400",-0.00858718682793502,-0.014551168722522,-0.00904992960961082,-0.00425763898236642,0.00787563556246207,0.00191592640017491,-0.00404105796711873,-0.00869335661975912,0.00320201923284325,-0.0059150056241617
"1401",0.000224205389453225,0.00691168773141393,0,0.00481047774018739,0.00257883570377193,0.000546270248383607,-0.00015605433203647,0.0112362353833357,0.0140046504949283,0.00743779921520837
"1402",0.0164969818071601,0.039001532955854,0.0148404084932059,0.0226063026798382,-0.00915557405220546,-0.00309439714888082,0.00811611269169399,0.018156915649902,0.00706626847904257,0.00184567420582926
"1403",0.0184330644862081,0.0252252896308165,0.0179977431019347,0.0280881839021998,-0.0188623301031637,-0.00721235988483604,0.0113019744346559,0.0159703275494441,0.00491158372363132,0.0103168479898337
"1404",0,0.000292921742659713,-0.00552501877991773,-0.00581835466358038,0.00747261124062959,0.00321873457347799,0.00275549029567945,-0.00314404757312581,-0.000698235399820168,0.00583515216558039
"1405",-0.00699460486229897,-0.00732060985955085,-0.00111091188872348,-0.00458002932519108,0.00200826359535,0.00174161950110441,-0.00106843302717075,-0.00210244346998434,-0.00597083174614632,-0.0119652153326775
"1406",-0.000871305053621985,0.00147497755845039,-0.00333703580461586,0.00178933100786272,-0.00499892224561871,-0.00364749091851513,-0.00290401909366345,0.00237005764408815,-0.0086267873785294,0.00146794543273732
"1407",-0.00690455926663291,-0.0191459584690391,-0.00446439347680483,-0.0117375144578268,0.00566825870104948,0.00239159013236745,0.00107293691398258,-0.00236445375239813,-0.00651021017474662,-0.00842810650609738
"1408",0.0198332995784838,0.0441441641539726,0.0112108294768711,0.03098363004042,-0.016137155863774,-0.00523021935965529,0.00734982337365486,0.0265999554696617,0.00921298873635923,0.0169993723911357
"1409",0.00193765303483229,0.00603958039920172,0.0099776868493977,0.00626121259229673,0.000391758825488475,0.000645321603136351,-0.00288796556534621,-0.00307832649310436,0.00482160067846471,0.00581391130596076
"1410",0.00501341308695147,0.00857634695033704,0.0120748212746327,0.00273738760263686,-0.0128654636537505,-0.00525409284682965,-0.0103659351966866,0.00385957541474014,-0.000127984642457113,0.00758667603917651
"1411",0.00121140460246449,0.000283596618301907,-0.00216938686191614,0.00198529434522365,-0.00532430522514049,-0.00139067558330164,-0.00600745297710059,-0.00589559637273285,0.00127973509905122,0.00286844636302375
"1412",0.000854629526162887,-0.00113360999869283,0.00217410333312351,0.0042114078973805,-0.000719398394960602,-0.000742334016893276,-0.00294429361658233,-0.00567322469499376,0.00325926005263955,0.00822316790061595
"1413",0.00163556462149161,0.000567465778748666,0.00108464773335926,0.00468676977792315,0.00503705924928788,0.00287949304355561,0.00217589033027155,0.00207471495896083,0.00121019169341396,-0.00531922193021361
"1414",-0.000497207686578793,-0.00255179765900493,-0.00216682336640328,-0.00883908932222821,-0.00167030144296076,-0.000648807068133195,-0.000310400673029232,-0.000776294577644054,-0.00757086176992006,-0.00784314027661215
"1415",0.000141980536476183,0.00454812729238929,-0.0010860388260252,-0.000247229342661193,-0.013546952210456,-0.00491074108707912,-0.000465237245993788,0.000776897679099608,-0.00551317374468951,0.00107795869947758
"1416",0.00113652992719193,-0.00226390750050254,-0.00543472403506051,-0.00148683255435178,-0.0140561325076567,-0.00502841572162416,0.00279371913252358,0.000776372983317675,0.00322310309988061,0.00861456835818042
"1417",0.00737852723387245,0.0116279990029442,0.0131148268680399,0.00918106207228031,-0.00852104204188386,-0.00243328348397853,0.0072744505701392,0.00517193521413728,0.0059756664532653,0.00391453712345635
"1418",0.00133784329314435,0.000841106885306919,0.00755149149820133,-0.00491754223549656,0.00487527158889112,0.00121994069049647,-0.000460722762815835,-0.00154348026702211,0.00102199158178307,0.00141799052216385
"1419",0.0000705658095359052,-0.00224080154889827,-0.00214151424716424,-0.000494225092292133,0.00205595958048388,0.000561926207879759,-0.000768698090699793,-0.00206138922817756,0.00344559722150595,0.00460174330616092
"1420",-0.00302411075000375,0.00842211155264549,0,-0.00148332116548333,0.00443207719176053,0.00084287133135863,0,0.00180762719567418,0.00998351169984457,0.00916132853008333
"1421",0.000423461753575882,-0.00250544909827033,-0.0010729797408694,0.000495320522999831,0.0165044244830836,0.00776682076104462,-0.000923134984927132,0.00180381899906323,0.0107661712426346,0.00523746664346136
"1422",-0.00817956317630764,-0.00586100735454365,0,-0.00915606924300294,0.00417974026717993,0.00176410472956179,-0.00261812032121045,-0.00565946661661765,0.00840915696314992,-0.00486276892515303
"1423",0.0060429886744926,-0.00364958860579034,-0.00107416243358638,0.000249707543371391,-0.000960856867708637,-0.00046356571771089,0.00385994231561382,0.00129347599834428,0.000494175060190116,-0.00453753155768599
"1424",0.000212071874894582,0.00338093405226769,-0.00322580148273177,-0.0102371864436103,0.00584916292396409,0.00259640112266757,0.00215336074495398,-0.00310106806129273,-0.0037661295069078,-0.00455828677532077
"1425",-0.000989563523945303,0.000561971729843513,-0.0086301677809919,-0.00201808551968674,0.00239001946422945,0.000369438366409902,0.00398997773454779,0.000518674928086327,0.00173523796643993,0.00070453633450196
"1426",0.000778306798012718,-0.00336823846738832,0.00326465790504038,-0.00480299095426884,-0.0043707165982162,-0.000647059802667438,0.000306022431082464,0.00259069594186578,-0.00649593545221427,0.00175991964506861
"1427",-0.00720814732678499,-0.0121089583710829,-0.0184382193754041,-0.0116841781229238,0.00518777120715241,0.00185057587402304,-0.00106988224162652,-0.0108528379473722,-0.000435842840422085,0.0010540966616186
"1428",0.00476913961519942,0.00940707891681702,0.00110514652774274,0.00950928391907224,0.014133709528743,0.00646401441049771,0.00397730359071335,0.00783682164137578,0.0230500679529013,0.0105300477460186
"1429",-0.000920961391475572,-0.000565006129355838,-0.0132451961353797,-0.00560075601580812,-0.00100434955778406,-0.00228760592368482,0.00502835287971792,-0.00596138498534637,0.00158321153584695,0.000347338084005111
"1430",-0.000850793465654975,0.000565325541751927,-0.0123042731220868,-0.00512032580414223,-0.00471249290167697,-0.000368713900468221,-0.000606486594225353,0.00286831923492104,-0.00103354817688583,-0.00486111622344032
"1431",0.0202964740117924,0.0293700668100656,0.0135898538829304,0.0221306659773308,-0.0166510048633036,-0.0068171513904316,0.00788842054955774,0.0176808286438026,0.00352991909841038,-0.000348877680432791
"1432",0.00389510274884008,0.0145405662438334,0.0134079911592158,0.0231621750609929,-0.00465460043874932,0.0012986454349746,0.00180633508814254,0.0107303683403202,0.0215295228426802,0.0111692034417417
"1433",-0.00568108502871634,-0.00919434471770775,0,-0.0127950568637192,0.00241890002205647,0.000463319752052715,-0.00646045058225897,-0.0123861518080045,-0.00682741027276867,0.00138079096165633
"1434",0.00278723497112665,0.0136462928451795,0.00441003331665257,0.0119638193076583,-0.00627358301750602,-0.00185159642877908,0.00393145201861134,0.0104942477820351,0.00364636873408197,0.00206822407648244
"1435",0.00333500206902415,0.0037696523206705,0.0109771999454502,0.00443349335475829,-0.0124642497278756,-0.00491634373339089,0.00376567345135759,0.0053189026008047,0.000119142350892609,0.00515995919531664
"1436",0.0152369529368044,0.0160944503816272,0.0162863736468242,0.026974128977066,-0.00393415451157741,0.00288953163695949,0.012154955594285,0.0191484303525737,0.0201881850903787,0.00684463933566049
"1437",0.00443391529664416,0.011615575566891,0.0106838856587941,0.0116999208340451,-0.0265781572495893,-0.00938855037296282,0.00518916706277328,0.00321399213031803,0.00286034093585119,0.0105370807807292
"1438",-0.00339567676114361,-0.00443644784117492,-0.0095137274768935,-0.0108568828963128,0.0120041433570666,0.00206441293839532,-0.00472006035712091,-0.00936423196287228,-0.00814906272149485,-0.02758157108499
"1439",-0.000818228637046392,-0.00786367926625975,0.00213465826896719,0.000477664959672497,0.00501141202797317,0.00252892384514958,-0.00859496802565829,-0.00273643235239285,0.00774652022581646,-0.00726389441688557
"1440",0.0005462194695669,0.00660498939033194,0.00212978216083837,0,0.00656561273564749,0.00233476462408588,-0.00463386337923688,0.000498987666397221,0.000116491962983467,-0.0146341610358031
"1441",0.0000682720326232733,-0.00839878984105313,-0.0106269955429268,-0.00596244821407399,0.00247713934166494,0.000558967607945604,-0.0117134451704872,-0.00299167748979456,-0.0015721671837613,0.005657667601356
"1442",-0.000418599780110274,0.00158800100323697,0.00537038978009718,0.00239907603438771,0.00115281577420978,0.00214218693643509,-0.000303883673175465,-0.00317918008828477,0.00285767771121659,0.0066807125953503
"1443",-0.00150770028585545,-0.00369991776292711,-0.00213636900395364,-0.000957457589125355,0.00781577106075426,0.00223057528067461,-0.00106412961491464,0.000759510169710875,-0.00529195140123473,-0.0104784481678606
"1444",-0.0106420691164141,-0.00822257580203967,0,-0.0148537444880531,0.0098773712467588,0.00370933003749485,-0.0146785559259105,-0.00758755286374002,-0.00163694238578882,0.0010589336079363
"1445",-0.00562140026178115,-0.0131049700395695,-0.0107068795419665,-0.00462046238611535,0.0107512675774553,0.00415704840419795,-0.000933955199065473,0.00331284943198051,-0.00562163130241533,-0.00705219856480976
"1446",0.00942147278918171,0.012195009321625,0.0119046927829405,0.0158805275572296,-0.00711826566460461,-0.00211560727964299,0.0054530754238149,0.00990603717974947,0.0148989931676462,0.0124289901219379
"1447",-0.00463217745637301,-0.0222220363557285,-0.0192513984914844,-0.00601244101019549,0.000564581949741072,0,-0.00232421056544629,-0.012826902706891,-0.00261110021146815,0.00596284678055925
"1448",0.0026398499575786,0.00930988342951045,-0.00327141045483359,0.00992005378515604,0.00371051368654474,0.00185527687001974,-0.00714531575765165,0.000764579657720921,0.00232703474505236,0.0013946092478001
"1449",0.00103889120541201,0.00623967422620186,-0.00437628913803645,0.00143767552585006,-0.00136624812131869,-0.000645129499976749,0.0084483644156792,0.00229091633098522,-0.00110271639514203,-0.00522287761086537
"1450",0.00408304091038447,-0.00269617181753401,-0.00439549436054276,-0.00669862949893318,0.000321990279935402,0.00101409626386983,0.00294766395963975,0.00101615439902836,0.00180126664260527,-0.0171508047357199
"1451",0.00716807345348935,0.0121654735127235,0.0121409595774455,0.0103563847329904,-0.0124710009997675,-0.00396071803639197,-0.00371231293520102,0.00888085845733255,0.00696013556150743,0.0217237170535389
"1452",0.0000685404368088172,0.00213692549205846,0,0,-0.0129539290667477,-0.00453120147894837,0.00434714578021,-0.000754508139878207,-0.00570247102296839,-0.00522833851815707
"1453",-0.00342146418897427,-0.00799614432709117,-0.00545262643871236,-0.00882005940818342,0.00841907772501638,0.00325119139980612,-0.00417397229750727,-0.00402688033317888,-0.00330200449837803,-0.00280311720481063
"1454",-0.0098875091374705,-0.0163887503014339,-0.0164471613374949,-0.00745533744789451,-0.0018007704646622,-0.00203698156682763,-0.00434632778152177,-0.0065707447810357,-0.00616098797743125,0.00737878512213519
"1455",-0.00638015143413428,-0.00273152165466517,-0.00780373644183474,-0.00605760248081522,0.00705195536815451,0.00241225070170126,0.00124733223170481,-0.000254178029882257,-0.000877296892294877,-0.00174399536590708
"1456",0.000558767824717865,0.00986018191029481,0.00561772646302994,0.00926365190811218,0.00692149719922019,0.000925722141349894,0.000155569923908194,0.00610682829291709,0.0028097109063383,0.0115304929006563
"1457",-0.00327859893563376,-0.000270964773239957,0.0011175575162059,-0.00314004297867065,0.0025068895410163,0.0000929575250852022,-0.00435918445454941,0.00126433267293535,-0.00735471018279843,-0.0138169849865292
"1458",0.00832769738199057,0.009223841487499,0.00669638644608028,0.00581533714859672,-0.00225881724992139,0.000276903323283006,0.00672387055271662,0.0101037095590799,-0.0100552276849962,-0.00490368285955811
"1459",0.0101334699995956,0.0185485700841777,0.0144123215999725,0.0103588792196971,-0.0138244871877187,-0.00471440097956055,0.00465995090436855,0.00975245193859453,0.00635575860923931,0.000704040312520915
"1460",0.00453483347957029,0.0102928546184431,0.00546442165878713,0.00786855354947869,-0.00926374152657738,-0.0063164003613766,0.00154609164827413,0.00990562858018107,0.000708269398043582,0.000351663888966014
"1461",-0.00259940081832033,-0.00548585873404117,0.00652160777947275,-0.00283918650693982,-0.00612329441344184,-0.0017759071666914,0.00941635230250548,-0.00662094611326314,-0.00442373499449178,-0.000351540264949435
"1462",-0.0166638997638006,-0.013396387238898,-0.012958703974295,-0.0154213007679753,0.0135704265624421,0.00421386509609056,-0.00932851174941496,-0.00987369546260097,-0.0107825823536826,-0.0151249139891453
"1463",0.000139197541015434,0.00559098596475827,0.0142231932353092,0.00963892286693135,-0.00640678261945904,-0.00335745672574961,-0.00355039232667775,0.00772808611939801,0.00365335686857904,-0.00464283041474622
"1464",-0.0138761103504662,-0.0238284818497299,-0.0204964250118485,-0.0205251170385472,0.0143016771687423,0.00477204840106316,-0.010069967568044,-0.0113800965316506,-0.0128297468333961,-0.0121995151716672
"1465",-0.00282852831168345,-0.00135582855575545,0.00220292894394114,0.000974606987582449,-0.00986155692169766,-0.00214188501170676,0.000625977440892767,0.00400381463821953,-0.00344551788743641,-0.00290588105193434
"1466",0.00290688305102105,0.00624662028871392,0.00769209969754869,0.0109541972064777,-0.00510413071516413,-0.00363905530588893,-0.0043788933629717,0.00822556573475164,0.00703629135608219,0.00255005608008707
"1467",-0.000565139828061945,-0.00026994820593762,-0.00545262643871236,-0.00770528873184073,0.0147276926530948,0.00636880349691382,-0.00581220302321339,-0.000494548717614118,-0.000542169605055598,0.00218020271517072
"1468",0,0.00242982318351803,-0.00657856886344477,-0.00145573721035874,0.00587108265302949,0.00409468324881823,0.0112183145395002,0.00766766400244201,0.00542402843348522,-0.000725227892248381
"1469",0.0104705120466311,0.0115807678244608,0.00993350956308503,0.016281913171325,-0.00818768289472005,-0.00199551413602173,0.00109347909074176,0.0108001919889995,-0.00455550554989503,0.00181427353995822
"1470",-0.00889184609889515,-0.0122472018524079,-0.00765040520925264,-0.00526069768071835,-0.000735530742777102,0.000837227695370313,0.00671152683616727,-0.0111703937042323,-0.0208948085369804,-0.017022771955908
"1471",0.00204861320960736,-0.00377355036769988,0,0.0048077188192881,0.00564384758095571,0.00241604162664233,-0.00744191375662495,-0.000982096574132507,0.00387447710180266,0.00847457402154794
"1472",0.00782540333832604,0.0113637324119289,0.00220292894394114,0.00789490681541194,-0.00943498077581229,-0.00454236270543384,0.00218666919119448,0.00958681093619962,0.0188078605356334,0.0179027562684033
"1473",-0.0226639853020209,-0.0160514937927543,-0.0120879335929149,-0.0163783420811374,0.0181461868996351,0.00838052770527353,-0.00498736109608111,-0.01266137682365,0.00114252553561278,-0.0186646826118815
"1474",-0.0120241994081509,-0.010875385876179,-0.00444962061386045,-0.0125481648883712,0.0148391383450324,0.00443287583599861,-0.010181734611507,-0.00838459558731108,0.00900954985255731,0.0014629624526632
"1475",0.000869551139677904,-0.00329873246686074,0,0.0019551603376371,0.00111225434674878,0.0000916396512218309,-0.00332334908525644,-0.00174084087061088,-0.00101195306232649,0.00803510311144295
"1476",0.000796175120991949,0.00193097827878441,-0.0100558207566921,0.00365862868250111,0.0016665423468909,0.000643528290911188,-0.00158782508033029,0.000248996998795104,-0.00220480267290191,-0.00471015522293972
"1477",-0.00347152668405337,-0.00330337353376975,0.00112875111443711,-0.00899161522824621,0.00332870126696516,0.00119442347000809,-0.00318084825883758,-0.00423410152427728,-0.00209012246205054,-0.00182014263204167
"1478",-0.0134987770925862,-0.00938935133316776,-0.0124015031779604,-0.0154485906398831,0.000947543958058628,0.000275193401452878,-0.0194636737620193,-0.0120059975910946,0.000239335718515754,0.00291761361802267
"1479",-0.00169202892339826,-0.00111531427008815,0.0159820129086623,0.0034867378848018,-0.00197251269685272,-0.000458649371007813,-0.0043930100161147,0.0075948952348488,-0.00628217665598985,-0.00400002006035627
"1480",0.0049374844723864,-0.00558183299659643,0.0179776462464949,0.00297848169028536,-0.000869784581451705,0.000641988901980195,0.0114397857818036,-0.00175900071828972,-0.00126432057954895,0.00438110108307055
"1481",0.0202388575130072,0.0224529708755306,0.0143484095918061,0.0175698748745647,-0.00561840127064284,-0.00201743195911919,0.00937128275019861,0.0148502927121781,0.0119965634194428,0.0189023340870691
"1482",0.000431465407974674,0.00329383164439445,-0.0021762246516942,-0.00194553614549198,-0.0100271975737898,-0.00413565439853247,0.00624311770656383,-0.00247978571553331,-0.00285933171082775,-0.00677854216455243
"1483",0.00186782174143163,0.00355665906878988,0.00109068456989947,-0.00194912798043057,-0.00056256983169467,-0.00147666715213868,-0.000636650591853138,0.00124291917576125,0.00101558636128574,0.00431032299677248
"1484",0.013625049398597,0.0239914417557368,0.0119823783531987,0.0163572086279857,-0.000964842447000902,-0.00055372583031299,0.00811876485995344,0.0144029247206121,0.0122344415401581,0.00357656282013474
"1485",-0.00212244900108005,-0.00213006535270888,0,0,0.00474981139721531,0.00166378263742795,0.00142106293915623,-0.00195860381134971,-0.00106130534130477,-0.0014254239409307
"1486",-0.00510434443638552,-0.00586967295338525,-0.00538198268502588,-0.00840731850671195,0.00392624974125733,0.00230801477866138,-0.00536128820541282,-0.00220711815675612,-0.00424946012952976,-0.00142760560061006
"1487",0.0080524040619534,0.00939338091955255,0.00108217847308434,0.00557172198130118,-0.00143668693834342,0.00128986468252701,-0.00174345826652245,0.00540787460149827,-0.0128030579715404,-0.00321664961115631
"1488",0.00466537980951243,0.00904003758986271,0.0118918237073187,0.00722715733181389,0.000159704413449369,0.00101160494421193,0.00651096569723553,0.00831284403673105,0.00378258774333373,0.00681249553246777
"1489",0.00021110399140678,0.000790606582562026,-0.00320488360930238,-0.000478272694444559,-0.00271752452766683,-0.000184085243632892,0.00394449921897966,0.00193971780819324,-0.00675912218754549,0.000712314306763551
"1490",-0.0049241884943414,0.00368605173756364,-0.00428749926353489,-0.000478642300978049,0.0009241687950865,-0.00039581587034887,0.00282876748647665,0.000484354003113197,0.000481794631464139,0.00249106907856311
"1491",-0.00141428065973115,0.00524680581856107,0.00107656585590643,0.00287286292358679,0.00577525779739596,0.00174930487436908,-0.00125361661563184,0.00217683088245257,-0.0102931857493174,-0.00887467772603245
"1492",0.00176998623138269,0.00182688257581409,0,0.0107421850317444,-0.000478252334617735,0.000827310948033233,-0.00266756271058288,-0.000482850525690637,-0.00182461381613697,-0.00107455759836994
"1493",0.00339234873891314,-0.000260782997411724,0.00537628546621538,0.00755807508062456,0.0021541111059411,0.00055082737529033,0.00881041626604917,-0.000241215581504028,0.00231540952703546,-0.00896381185338879
"1494",0.0030285534927601,-0.00286598318636921,0.00320855139450216,0.00304729909870494,-0.00923615150062107,-0.00284491549716193,0.00405495503338038,0.00942023067412601,0.00401218237082057,-0.00108533151390944
"1495",0.000421470678664271,0.001306551927994,-0.00319828951820844,0.00560887346468997,0.00442033034096423,0.000920472454073673,0,0.000239201771688347,0.00387502412509044,-0.00217317058423616
"1496",0.00680818359000912,0.00887267012537873,-0.00106920670276123,0.00511284958355507,-0.00760148404405658,-0.00193054946343452,0.00124268242664161,0.00311024428089612,-0.000904758729105781,-0.00181478263702284
"1497",0.000488318732732251,0.00439730313135134,0.00428233680047385,0.00300564689299843,-0.0116098626486748,-0.0042390795314996,-0.000620683248861331,-0.0007156031053559,0.000724479350117102,0.00472724539946046
"1498",-0.00613234801281781,-0.00283305513795251,-0.00426407658837935,-0.00437985488583226,0.000733852934111878,-0.00194251818285007,-0.00667473311138933,-0.00548934736449225,-0.0084454905363941,-0.00904819863907314
"1499",-0.00371563907356753,0.00490713267594711,0.00535325932910813,0.00439912240358509,0.00749938325997102,0.00222495626734243,-0.00125033897947679,0.00551964662213034,-0.00146005966599916,0.0062089023060381
"1500",0.0117521428190941,0.00429222289462694,0.00958440859941656,0.00253564979558218,-0.0149676005152212,-0.00527253064287847,0.00625877405264941,0.00811462664866491,0.00188872838942511,-0.000725868225068038
"1501",0.0111285496038149,0.00875380880817045,0.0150336084790705,0.00698611584337216,-0.0101848905636908,-0.00390518555510788,0.0102628202883912,0.00639202450162912,-0.0143517390616426,0.00254264592044251
"1502",-0.00742875318575975,0.000765777852314908,0.0157565204699701,-0.000459266719449514,0.00331917516995528,0.00140009567560573,-0.00140238692086336,-0.00352849153163792,-0.00240621912134487,0.00362325082674775
"1503",0.00575196444593273,0.00586565731992406,0.0134434936708701,0.00597562937794849,0.000165457751373443,0.000652667026409537,0.0113904361228794,0.0144002100525367,-0.0121219987368173,-0.00469318791637974
"1504",-0.00907728900232796,-0.00938105721731675,-0.00612254458206762,-0.0114233045810979,0.0109155445305977,0.00270121533982848,-0.00308545412852035,-0.00667207543768067,0.00375637647921812,-0.00181354069069395
"1505",-0.00308096880824116,-0.00204776047126831,0,-0.00208021258882496,-0.00179961036078979,-0.00102144354104827,0.00139267556983302,-0.000486998871302324,0.00180872573057145,-0.00327037887043391
"1506",-0.00421509418821397,0.00102591824609122,-0.00102678625943819,0.00301074426711812,0.0035967989960819,0.00205789371165999,-0.00494519986319453,-0.000973768465308944,0.000996164892173024,0.0102077748250822
"1507",-0.00134050588403822,0.00435567610913234,0.00102784163310399,0.00563566224019363,0.00335551244438448,0.00204534053212235,0.00124244410019303,0.00316869529696806,0.0023635091576284,0
"1508",-0.0108080281078219,-0.0142856914755879,-0.00718661934418729,0.00367454526270738,0.00570918039420176,0.00231869036328303,-0.00604939640719948,-0.00753190369110734,-0.00384717662330147,-0.00288700503424477
"1509",0.0169963968496489,0.0170807097329388,0.00827285949570933,0.0148742261335719,-0.0172737405110055,-0.00527494758029079,0.00920740232890527,0.0122399575136123,0.00921895517959803,0.00542888193349578
"1510",0.0256302654981806,0.0145039148175474,0.0246153130532256,0.0196168934855425,-0.0133684947806785,-0.00455862874218582,0.0162362118694279,0.0133011128273477,0.00709785194178858,0.00359966281133017
"1511",-0.00225972414376852,-0.0135440953261109,-0.00900881654300201,-0.00707675688843867,-0.0135494916592457,-0.00514048687159696,0,-0.0152742481168189,-0.0120733040641454,-0.00824960277536924
"1512",0.00439174515400143,0.00711918917394971,-0.0040405414994803,0.00200472435241905,0.00390002601197526,0.000469909408553182,0.00608620210438837,-0.00169689487259683,-0.00471460926888234,-0.00433994176907604
"1513",-0.00273269976590762,-0.000757154821817263,-0.00912770626654535,-0.00755717985219717,0.000422352106863366,0.000563367268517245,0.00151254430567449,0.00315614132396935,-0.00629524424962291,0.00181617565745906
"1514",-0.00287729099798184,-0.00202137428893745,-0.0133060940934759,-0.00895868254896315,0.00658536109721863,0.00243976489438213,-0.00196305097175398,-0.00847047776660925,0.00708778178269132,0.00253807371799342
"1515",0.00254196581243704,0.00101267211899536,0.0134855338761326,0.00429381099322446,-0.000922695887488612,0.00056192732383642,0.00378253093609948,0.00488160756672995,-0.000435930498703718,-0.00144667207169502
"1516",0.00794992765952585,0.0174507900756165,0.00818838309982328,0.00877572496154255,-0.00277041109964615,-0.00290015600373894,0.0024118476290298,0.00777283982169985,0.00928401117564914,0.00362186399421871
"1517",-0.0000679713918859681,0.00422563002204646,0.00304550678002458,-0.00803016629054754,0.00892333911414478,0.00319041363576433,-0.000150301415831056,-0.00385640955040167,-0.00567970133793549,-0.004330618978589
"1518",-0.000680089836984865,-0.000742592003032949,0.00607296969320581,0.0042723583569011,-0.00275361741505298,-0.000374245272929397,0.00150414685122158,0.00435512525601256,0.00298022479796622,0.00652420086718264
"1519",0.000680552673941959,-0.00346783238967197,-0.00301826750774081,-0.00425418296276836,0.00460182255130936,0.00243252572411778,0.00465532860069207,-0.00192727598128251,0.00631425680450537,-0.00432122496650611
"1520",-0.000136438745114931,-0.00472273245937682,-0.0121088349302643,-0.000899562843790891,0.00208209733116016,0.00130709397833728,-0.00104650474136181,-0.000483002313073522,0.000553617132795337,0.00108497613651792
"1521",0.00646054952071085,0.0107389534694291,0.00408571415919545,0.00562700103852531,-0.00997322356685204,-0.00456806363243523,0.00224460446328223,-0.00217314714442074,0.00430379358021993,0.00433527532181133
"1522",0.00222998692458276,-0.00222374099229328,0.00406931518557041,0.00223786591463648,0.00772331183136199,0.00280984836628462,0.00597171094195192,0.000967876707268722,-0.00159173547872404,0.00647484275670118
"1523",0.00539306231058156,0.000247278417748742,-0.0101317195621293,-0.00156319367649349,0.00191562268032253,0.000840301513144182,0.00504634730470443,-0.003384712242673,0.00355633094748486,0.00285914600816461
"1524",0.00160954731494334,0.00049540691187433,-0.0081883830998235,-0.00536775165805048,-0.00149655611169752,0.000466838082797016,0.000147651705014296,-0.00388156525620575,-0.00281047843600513,0.00106912297437733
"1525",0.000267964647804764,0.00569171622332143,0.0113518950970086,-0.00359801480028232,-0.00349735880856072,-0.00167898766650076,0.00118088444847131,0.00487115354979051,-0.0109675199021344,-0.000711914167553562
"1526",0.00562184777409258,0.0135335372770813,0.00714293087019024,-0.00338529127439413,-0.013704227008033,-0.0066332338620797,0.00412941897417052,0.00581636893852511,-0.00477018962669051,-0.00213755737961818
"1527",-0.00119807158378205,-0.00194209655551891,-0.015197579343194,-0.00701985172689479,-0.00364335851855002,-0.00206884181264966,0.00102800338109654,-0.00578273442165522,-0.00224090266694921,-0.000357010471621177
"1528",0.00393145790411875,0.00510815863461445,0.01337454112965,0.0111744538031255,-0.00552709779214411,-0.0015081049164134,0.00190731215550044,0.00290792174323418,0.0043671597140813,0.00571428109331551
"1529",-0.00391606207093687,-0.00121019564210767,0.0101520654363589,-0.00473601123534928,-0.00171021007052508,0.00056645458242377,-0.00922524132891223,0.00338360019923245,0.00745386025672823,0.0113635906775538
"1530",-0.00246534985210822,-0.00411911548823396,0.00201023079447005,0.00203919976401834,0.00488254071487959,0.000849043535311234,-0.00576427815787017,0.00120389607839844,-0.00610398290765168,-0.000351118811761197
"1531",0.0102873026638322,0.0104623479157988,-0.00300907382538362,0.0065580555979099,-0.0129846587436601,-0.00339732534120452,0.0066895732585095,0.00384923276806948,0.00155086851521458,0.00386373583612265
"1532",-0.0112403404207178,-0.0276908848554497,0.00100590278740764,-0.0132554622744313,0.0128090309356581,0.0057764794326205,-0.00206729805624628,-0.0134197376179883,0.00340664608374075,-0.00349897458315218
"1533",0.0100973238348474,0.00693391660565768,-0.00301501104152291,0.00113865487922071,-0.00888718332272964,-0.00357783559957037,-0.00133221941389206,0.00607251575151024,-0.000246870370370411,0.00386237920578703
"1534",0.000728355361654387,-0.00270525568342606,0.0131048943980894,-0.00113735981891339,0.00819120960407527,0.00302350927003858,0.00177832550724721,0.000482490770405519,0.00265492702775694,-0.00139907150236718
"1535",-0.00132267426662325,-0.0120839150527655,0.00298512118005911,-0.00887954917336542,-0.0022234640023161,0.000470950901004352,-0.00473293018350296,-0.00627367998111006,-0.0033869265557418,-0.00385290912519543
"1536",0.00556401653759742,0.00848743244706318,-0.00396827891161644,0.00735120812372547,0.0038568787119091,0.000753571214204607,0.00995675779086369,0.0106848026051283,-0.00166824645744557,0.0038678114512305
"1537",-0.000197878010279151,-0.00594085753655715,0.0109560506889923,-0.000455981011356577,-0.000768895309459006,-0.00103506003675646,0.00103012425924498,-0.00336401811909404,-0.0115739921952223,-0.00350257911454177
"1538",0.00164725329463011,0.00821742169921524,-0.00689640444479245,0.00273777422747767,-0.00247748811006143,-0.00103605677044161,0.0058796760129689,0.00168761677868723,0.00118974329097821,0.00175744514794096
"1539",0.000855240812945413,0.00493940709049845,-0.00396827891161644,0.00500562847949992,-0.00813835665335017,-0.00348887711012058,-0.000438378430371422,0.00553530180241157,-0.00525358687381061,0.000350872390607826
"1540",0.000920277145950443,-0.00737311616119007,-0.00996016686119339,-0.000452677556651682,0.00906847154333978,0.00425772359536514,-0.00394753860631181,-0.00526523172381677,-0.00440111277457822,-0.00140306948977265
"1541",-0.00118203028308284,-0.00321841294767111,-0.00301826750774081,-0.00362390778320731,-0.00290974426280488,-0.000942152994297119,0.00117452879616464,-0.00433150949715189,-0.0163562418810391,-0.00421490567380778
"1542",0.00749443889257817,0.011177677044004,0.0151362399562276,0.00204571599275849,-0.00497845660847396,-0.00160321493019877,0.00689021992707484,0.0113582113220254,-0.00276061256935711,-0.00388012635360513
"1543",-0.0124631872303997,-0.0132649894585879,0.00298204376072975,-0.00884752896143393,0.00301921380582915,0.00217283528137635,-0.00844489902996171,-0.0074073449862484,-0.025043455545697,-0.0113313996413342
"1544",-0.00607911602637501,-0.0164301716558926,-0.0118927104598939,-0.0137331651097351,0.00584801675050817,0.00197857702189408,-0.00778256808907474,-0.00698096947575555,0.00779181843909371,-0.0114613456196369
"1545",0.00977309706777696,0.0151863647846833,0.0160480220933741,0.00440926662168128,0.000684077626547097,0.00122344470659885,0.0085839939295238,0.00509076284602972,0.00229331680950451,0
"1546",-0.0190270323618447,-0.0309152515073503,-0.0138203691086599,-0.0134008727423505,0.0196532442709683,0.00770348533255705,-0.016874940609535,-0.0159188267601392,0.00895597170062135,-0.00471015522293972
"1547",0.00684533104438367,0.00694639851315082,0.0190193637704128,0.00562064342987401,-0.00578204612088351,-0.00186437351401447,0.00880598742512095,0.0137250960746098,0.0121809320249042,-0.00182014263204167
"1548",0.0125985922174356,0.016607114810312,-0.000982488039925733,0.0109451854357145,-0.00295015655702369,-0.000466947881735402,0.00769341373843679,0.0108803382944003,-0.0105619894343746,-0.00619988201925725
"1549",-0.00197508974462657,-0.00276465169163975,0.00393316128781218,-0.0046072943769665,0.00185989459168723,0.00140173419850309,0.000146883252080121,-0.000717797612738713,-0.0101572551523531,-0.00440368522061918
"1550",0.00329797536182608,-0.00453621371646051,0.00979410816240267,0.00231462100042434,0.00544590878435813,0.00249454177308439,0.00190837451171566,0.00694131895784378,-0.00366011764705887,-0.0070032599178137
"1551",0.00532494911573522,0.00405043991411436,0.00581968402624078,-0.00946678965171266,-0.00529867594798783,-0.00233000646633619,0.00747274114444263,0.00499167561632397,-0.000918387550270405,-0.00371197812652269
"1552",0.00895896273887975,0.0115986719689709,0.00192870615363683,0.0121211477166445,-0.00287475104967405,-0.00102787620588485,0.00770801696781231,0.00402091386618753,0.000525292176126957,0.00931452061308158
"1553",0.0013611534643434,0,0.0125120826956542,0.00483657560658313,-0.00907303810037541,-0.00317894927788676,-0.00375245153988213,0.00235558683747761,0.00557810061759745,-0.00553713659489818
"1554",0.00181255129053182,0.00672960536613765,-0.00950570985025778,0.00275040495042345,-0.00770165580643689,-0.00384607959148831,-0.0036217167974294,0.00164504255527298,-0.00352407501204921,0.0066815377053342
"1555",0.00426425676869102,-0.000742411498885542,0.00479857444511067,0.00868584664554395,-0.0104343821740989,-0.00508529783750222,0.000581542897830634,-0.00351932116714482,0.000131017091741237,0.0029498120940703
"1556",0.00379529407629731,0.00322104737512485,0.005730216404771,-0.0054387225026955,0.000958303488992174,0.000473281291103911,0.00392329496977251,-0.0014131154043906,0.00183352751728982,0.000735284073664522
"1557",-0.00224302635727458,-0.0027167345208724,-0.0104460165635155,-0.0113921471906177,0.00722621139748725,0.00274350935550305,-0.00361851506136923,-0.00589438748703286,0.00784363004628963,0.00220426929571249
"1558",0.00141316464707497,-0.00247673528298287,0.00575803330775204,-0.0094490145653966,-0.00103720282349007,-0.000849210407496637,0.000290670344416766,-0.000474261963672951,-0.00343730457957969,-0.00513193244750831
"1559",0.00532374842567829,0.0139031185629406,0.00572517424143593,0.00418795937202909,-0.00302845884180691,0.000283393776806529,0.00537316455484182,0.0163739514528531,0.000130085900557519,0.00736920964057641
"1560",-0.00132018371470755,-0.00171412666837434,0.00948777930195432,-0.00903612344957649,0.00468658187163506,0.00349240918360216,0.00043346409449696,0.0002812058801962,0.00208229447277497,0.00219455661418477
"1561",-0.00551876826660458,-0.0139809607855373,-0.00469914698676854,-0.0112229719545273,0.00760204279968324,0.00329310119015913,-0.00274351542695206,-0.00726533871885915,0.0089610714285715,-0.00583944890513199
"1562",-0.00232306668775006,-0.00248770313983138,0.00566549490551549,-0.00709373452615458,0.00677309830674755,0.00309395670665702,-0.0070941136496544,-0.00613795841109743,0.00450506485696156,-0.0073420437609536
"1563",0.00698519721050062,0.00573583974795877,0.00751178511096762,0.00571545970786991,-0.0111556433423118,-0.00383250482975772,0.00583259834438765,0.00356294678950975,-0.00454899404729647,0.00702653066856218
"1564",-0.0085428377407234,-0.0116540530493443,0,-0.0101822610077458,0.00964480388667655,0.00262740744674983,-0.00333441376413235,-0.00591679868127915,0.00566393144313371,-0.0044069196129316
"1565",0.00803332883045571,0.0102862899285232,0.0037277858553606,0.00382803662796194,0.000767712680703081,0.000374420140776044,0.00610907496461244,0.0128572118473131,-0.00447998080000001,0.00184431274578434
"1566",-0.00417734376694434,-0.015644742346657,-0.00928485269585322,-0.000953680034038618,-0.000937856278441007,0.000748484879153244,-0.000670409586320919,-0.00188080851484451,-0.00199291542283031,0.000736442796368086
"1567",0.00800262767268767,0.00479342948696604,0.00937186912011834,0.0143133627543379,0.00119479398058364,0.00102831251520441,0.00744056402620585,0.00894982736543137,-0.00334967781017526,0.00919792752690629
"1568",0,-0.0100428800275294,0.00464252955882816,0.00376271981180798,0.00852076429867599,0.00429588620359378,0.00159323249222365,0.00396820903132156,0.00413650462683246,0.00510390617331535
"1569",0.00307322381356157,0.00710125916234405,-0.00184838933703724,0.0021087807114557,-0.00506903716212381,-0.0018600139761068,0.00462693372601586,0,-0.00585738925169044,-0.00943056091566707
"1570",-0.0039570476124936,-0.00528828197206366,-0.038888596698521,-0.0107552581588561,0.00753124589102128,0.00265880131152274,0.00316644469431981,-0.0179027354025906,0.00142441569616869,0
"1571",0.00493407343489571,0.0108859223444255,0.012523839624667,0.000472909381782127,-0.00405408462850521,-0.00195375561006839,0.00258254319534146,0.0187026275203781,-0.0144824790131568,-0.00476013385914431
"1572",-0.0101388874463728,-0.00500868112998132,-0.00380571166638954,-0.011811899256527,0.00898952001259468,0.00419513367825441,-0.00529479581822978,-0.00720415309926825,-0.0111526410684805,-0.0169242426921778
"1573",0.00405849411878423,0,0.0410693643582303,-0.00286898143013248,0.0119360054167732,0.0039917141896566,0.0146737459748032,0.0203649629256342,-0.00291914689628192,-0.0011226621444842
"1574",-0.00449153894710663,-0.00604058049055201,0.00550467379214181,-0.00239763608417642,0.020184451072824,0.00314430505253593,0.00269394092603581,0.0142232370587836,0.01676761672349,-0.000749411160418934
"1575",0.00676759841797692,0.000759455464496073,0.0100364844129619,0.00168239584720409,-0.00765355188071015,-0.00322654124208743,0.00933266530989108,0.00226191052217217,-0.00425360911267092,0.00299958406858414
"1576",0.00345660012377058,0.0055668319667328,-0.00812990741340436,0.0098369013342916,-0.00246157740637876,0.000370025952773689,0.000420609080254986,-0.00112846789049947,0.00775494196227822,0.00635520752959895
"1577",0.012248765164637,0.0158531475802917,0.0209468515373987,0.00950334703969058,-0.0137358657927876,-0.00415952602009495,0.00588133786773626,0.00610054590302456,-0.0168905443299999,-0.00222887210996559
"1578",0.00327733101026539,0.00569699035098603,0.0115969140572698,0.000941481901095775,0.00191781368999377,0.00111363226218875,0.00487250354754121,0.00381760824767863,0.00199006965174142,-0.00409532978060922
"1579",-0.00244988225230225,-0.000985114550059452,0.0017635572251713,-0.0152834125743566,0.0148998659423445,0.00556302956957255,0.0058189589322899,0.0123042306746488,-0.0470043419992517,-0.0123363959983461
"1580",-0.0231739042640957,-0.0219428256535333,-0.00792239125649141,-0.0243553508447762,0.00869365997648019,0.00221336619399248,-0.0249313330903618,-0.0227623812968403,-0.087808261642409,-0.0299015704037351
"1581",0.01476297788584,0.0143687635848639,0.00976041426970631,0.0205582060529563,-0.00821218614461483,-0.00285189279761011,0.0158217421602813,0.0174129261726217,0.0113472319145111,0.0105344659073492
"1582",-0.0146114910657665,-0.0280817048644068,-0.00702982427539389,-0.0158273732201655,0.00664015408405172,0.00184471063803282,-0.0120987049542109,-0.0111137312998252,0.000527048180864798,-0.0146718133830123
"1583",-0.00625403971758498,-0.000766834707973896,-0.00707959256708202,0,0.00244325691489022,0.000552694888491967,0,0.000449657979081586,0.0107624599519254,0.0105799947329301
"1584",0.00869371786878359,0.00690881861798753,0.0106950563067425,0.0146199599950394,-0.0021123160268689,-0.000552389585591451,0.0115429512458864,0.0146033217949166,0.00871182407940818,-0.00232653110253789
"1585",0.00443822159395713,0.00482850549839142,-0.000881815371229888,0.00480291173418368,0.000733276223188195,0.000552694888491967,0.00139156777853433,-0.00221400957784823,0.0179374989448771,0.00310924862864859
"1586",0.0103090026102353,0.0171978859224107,0.00970865285166234,0.00478017754410343,-0.00349840672520474,-0.000644512515162621,0.00583674818201319,0.00199733675653602,-0.00739658480333205,-0.00619922233375714
"1587",0.000633617609270276,0.00795607420717848,0.00611892080499388,0.00594656579798336,0.0025307204335201,0.000460816743149683,0.00317752511854708,0.00442950852057389,0.0108853736526382,0.0109162716021534
"1588",0.00405381530476756,0.0051802235921774,0.00521313342637408,0.00898571401799031,-0.00431581430073846,-0.00110483481990642,-0.00123975386839836,0.00308718530507934,0.0235600933569451,0.0131122044342977
"1589",-0.00176651457498866,0.00294455428672968,-0.00259304880379163,-0.0100772628228746,0.00915967778957172,0.0035947902856508,-0.00455009861868261,-0.00395681875531517,-0.00508367559543632,-0.00570989639238018
"1590",0.00669860371398046,0.0149254820445135,0.00606565534603631,0.0104165421344098,-0.00364669979605681,-0.000367792863536831,0.00775700096209797,0.0134626942500304,0.00986444511065376,0.0133996281898012
"1591",0.00238576934114487,0.000482181490012223,0.00775203632564092,0.0142925183818192,0.000569221643019313,-0.00018332207576377,0.00975928776517176,0.00413726509832957,0.00330288819459823,-0.00755569810693069
"1592",-0.00876752233775102,-0.00578294564381832,-0.0111108735937188,-0.0108569376836294,0.0102731550694575,0.0032657692498026,-0.00680618950617917,-0.00303605246743732,-0.011627113213501,-0.0178911993642445
"1593",0.0092874244134078,0.00484722654968994,0.00432125962797869,0.00794007478776471,-0.00129015704370306,0,0.00383739949659501,0.00478577272577385,0.00574018137807242,0.0127906433562244
"1594",0.0101404483160719,0.0125421727457831,0.0137694278328364,0.00834087869349442,-0.0235770166497653,-0.00852805339286211,0.000819375729631977,0.00974246389783273,0.00119784387257416,0.0110984797220384
"1595",0.00254058385291467,-0.00214401690562793,-0.00424455638892696,0.00137893382452581,-0.00248086490912514,-0.00129459120893516,0.00395642065202217,-0.00171522488946518,0.000422253513188808,0.00113548788016282
"1596",0.00506916519384903,0.00429701280147587,0.00170506451614361,0.00711316972837306,-0.00389619070198199,-0.00138964567002431,0.00584335917886536,-0.00536945736350702,-0.0124515587387221,-0.00340260002939397
"1597",0.00455107290604628,0.0125981290646164,0.00851057459203064,0.00774701058608529,0.00158157118476798,0.00120586151839208,0.00243174918023437,0.00539844407881751,0.0148169392072608,0.00455228966012333
"1598",-0.00281618091113744,-0.0103288083505114,-0.00759470445405763,-0.0072350752753555,-0.0025761700335053,-0.00018532469822985,-0.00512130336514716,-0.0124570557498128,-0.0115822611183781,-0.00037763835250948
"1599",0.00325378235659235,0.00403239387169751,0,-0.0077430545073407,-0.0107461307104891,-0.00565137333660626,0.000270850111090626,-0.00282732686696896,-0.00859308299968875,-0.00453344997004712
"1600",0.000795643721724471,-0.00496093626553207,0.0127549453075584,-0.00918085502054711,-0.00766353512854767,-0.00177024747602161,0.00148980904297624,-0.00937838770574895,-0.00838118158820145,-0.00455409573522136
"1601",0.0103336833674725,0.00189956504031086,0.00671708744400479,0.00463290790795456,-0.0108618534583176,-0.00401364209420141,0.00527395305963507,-0.00440346303366035,-0.00447876205556108,-0.00343117818564065
"1602",0.00538621674687922,0.00402801732317348,0.00917437018870526,0.000230635101201582,0.00669154489126877,0.00262412430273784,0.00887782182576125,-0.00309599701344876,-0.0230751980708975,-0.00229530155362823
"1603",-0.00469526565268563,-0.00330413992329148,-0.0148760807371786,-0.00345786652305935,0.0103972685619598,0.00476690400657898,-0.00319972380813327,-0.00155271019043024,-0.00401105979309735,-0.00115036996924256
"1604",0.00967710593384585,0.00710389208961182,0.0159395585119806,0.00439501432745959,-0.0126518109740063,-0.00539523216318727,0.00628662390752766,0.0135525241466681,-0.0225221052284915,0.0049904142640429
"1605",-0.0000598816619380438,0.00352726652571134,0.00660596921484147,0.00253355333439642,-0.00119612682916237,-0.000748455790238411,-0.000531391943199178,0.0054797798810875,0.0308994261364461,0.00649353610594772
"1606",0.00143764532389334,0.00234271858529711,0.00574256323812539,-0.0020677370795501,0.00786859481754543,0.00262085590901107,0.0046544892858027,-0.00893779495936309,-0.0165777833251103,-0.00569256107987448
"1607",-0.00741743448666643,-0.00864875471685123,-0.0106036337784639,-0.0110496599772396,-0.0148505350111573,-0.00793530778559803,-0.024755236995413,-0.0217775427452259,-0.00707407408661687,-0.00458016862487476
"1608",-0.00289283348808667,-0.00495146190448448,-0.042044535421634,-0.00744863725632317,0.00473784988732628,0.00103552810178176,-0.0139810929800924,-0.0179899050962512,0.0202364632372829,0.00460124309412979
"1609",-0.000846469751980883,-0.000711120831067835,-0.0180721184362259,-0.00867759072561247,0.00137174848664068,0.000375842488750777,-0.00385451917133384,-0.0137389519359189,-0.00631458282211894,-0.00381682028174757
"1610",0.00598900019204085,0.00497964200557832,-0.00613512950310957,0.00544148965442459,-0.025342665302083,-0.0117459577222248,-0.00995041182611756,0.00371459250146855,-0.00201846598454203,0.00919547400448573
"1611",-0.00649438918700229,-0.00542690974729476,-0.0167546880994722,-0.012705775531794,0.0112439054969367,0.00408882386258425,-0.0199606633426922,-0.0168862350183661,0.0100381822594133,-0.00645409096761351
"1612",0.00369219292958234,0.00711760744966727,-0.00538124942925544,0,-0.00243201722442865,0.0000948198890193819,-0.00954279602916697,-0.011529524018882,0.013869279628135,0
"1613",-0.0143521937469149,-0.0209659723929581,-0.022542849003957,-0.0181125381442067,-0.00339624270731576,-0.00274601659607854,-0.012223316964649,-0.0211854218277148,-0.0203364964228931,-0.0118455806241523
"1614",0.00550635788643428,0.00986520449778805,-0.0119925679918104,0.0148058512392708,0.00529887806365537,0.0014448744622515,0.0024750247979255,0.00437753713570577,0.0193398823079434,0.0123741931688792
"1615",-0.00480687342433372,-0.00381226957723713,0.0289449121700298,-0.0121983545614835,-0.00923489581471804,-0.00256338061356109,-0.0116179456002435,0.00750609930694734,-0.0093765954646764,0.0038197756843481
"1616",-0.014000856300339,-0.0150680557417878,-0.0381125107867263,-0.0179176329316113,0.0138052040885781,0.00485448751573325,-0.0107256463314803,-0.0206685446985225,0.00214455378672063,-0.00456618679793841
"1617",0.00905281093135701,0.00801355091707445,-0.000943271079539287,0.00838281431273891,-0.000606454237205289,0.00123149810130729,0.0187138272975125,0.00490838927432247,0.0074527373833313,0.00382265631848155
"1618",0.0127206000468476,0.00939525456786305,0.0387155622406703,-0.00513457418471241,-0.0178794397780715,-0.00775789933277327,-0.000583364864606195,0.0144075907554795,-0.0238042922713271,0.00228477333300514
"1619",0,-0.00167052808903945,0.0127272021740106,-0.0135166747598274,-0.00477158503638386,-0.00247903671840588,-0.00875286963831712,-0.0122773942143748,0.00495200333847534,-0.00379945755776012
"1620",-0.0103154428646587,-0.0098018793047745,-0.019748630928825,-0.0189335526231873,0.01189802474329,0.0024851976145448,-0.0153051853897871,-0.0216912629836181,-0.00515157525531462,-0.00877181068797406
"1621",-0.00827720782696717,-0.00120691858009259,0.00274749939992924,-0.00685633179777767,-0.0143029672624183,-0.0044814500038175,-0.014646396519102,-0.00747387768555774,0.00750469043151969,0.00115427429577508
"1622",0.0152086776193512,0.0120859058649017,0.0237439057184301,0.0212219123506452,0.0156682487543551,0.00756652470091645,0.0304870622065543,0.0256019778925185,-0.00379884543761644,0.00653342551185299
"1623",-0.00627275287224438,-0.00740368527575408,-0.0312218812198769,-0.0157735589559027,-0.00236690344977308,0.00133063162776859,0.00250175307496114,0.00244788748729663,0.00515917432484025,0.00420005822399827
"1624",0.0077219826193351,0.00986520449778805,0.026703539229709,0.00915757108137183,-0.00527108988074032,-0.0023731989279927,0.00132137791484688,0.00366189846207932,-0.00490953681742734,0.00228141593051934
"1625",0.00790566416488447,0.00333571760402052,0.0170401911879823,0.00428572262057569,0.000529798836262252,-0.000570909607881642,0.00161324192264289,0.00997344292743607,-0.0122598411524305,0.00189678735838483
"1626",-0.0138170110043331,-0.0189979760031916,-0.0123456112433225,-0.0308734411931526,-0.0103280987254335,-0.0137104408838633,-0.0300102505876776,-0.023603348662532,-0.0116552557460359,0.00151455709395831
"1627",-0.024778227226389,-0.0326797496301096,-0.0410716398285941,-0.0448072328281519,-0.0164130571290385,-0.00453700389701517,-0.0390887857029548,-0.0434137346223759,-0.0535262900230122,-0.0325141227318189
"1628",0.00321016443014943,-0.00900907154090702,0.0363129066936978,0.0143709942386452,-0.0169582289488038,-0.0105701485162695,0.0117795886052503,0.00489228120642604,0.0117314322286639,-0.00625247726745759
"1629",-0.0126358204840716,-0.0154040286334264,-0.0278525573515637,-0.0203152346324078,0.00415121418723463,-0.00245079318774599,-0.00636438860301569,-0.0190053808573135,-0.00895644120856198,-0.00432562145749138
"1630",0.00961399967864929,0.0118641450433667,0.0129390335611288,0.0212823164419464,-0.00891110894336289,-0.00117885189348188,0.0184346521970997,0.0177812029316697,-0.00371176470588241,0.000789878627295737
"1631",0.00990105099651672,0.00726355743720442,-0.00456194616802086,0.0157625207890999,0.00648866511092172,0.0040333154035157,0.0149570977641653,0.0104303292388304,-0.0420345181660766,-0.00276239324015415
"1632",0.00586982394462265,0.00463523708535574,0.0245787580794687,0.0200656674222264,0.0102230634778828,0.00538863853525084,0.0178491269799961,0.0198707497950887,-0.0197835392271182,-0.000395720742039196
"1633",-0.00409750703306977,-0.0066648439441952,0.00808614983939426,0.0057471354443428,0.00683720174906233,-0.00116937980880294,-0.0043466279009835,0.00961567287037712,0.0273417193834444,-0.00514652842086805
"1634",0.00585990058013985,0.0118708756515817,0.0124777078538023,0.00311707868244171,0.00201487931831301,0.000380703239706515,-0.00526846697187466,-0.0045114514525656,0.0169590796997812,0.00636692819458662
"1635",-0.000929638757096396,-0.0104564433424565,0.00704233465473769,-0.0178665818605667,-0.000634208029164141,0.000390743728601706,0.0116522649933863,0.00881163473711988,-0.00891599130477971,0.00395407799903147
"1636",0.000434083794563112,0.00128879696417683,0.000874235645459631,-0.00922736316653971,-0.00299023504958562,-0.00195239856904006,-0.00433815657600922,-0.00349383180352547,0.00574756337157267,0.00905876382185755
"1637",0.0107887564597449,0.00180169701962352,0.0131004129375549,-0.00638640697308734,-0.0340882383751223,-0.0168233287247755,-0.0105168195297473,0.00776345340478168,-0.0219480043390426,-0.00234196863799574
"1638",0.00570500656689465,0.0107913875215961,-0.00689636764254531,0.00133890384404833,0.00969326325925168,0.00587017342110063,0.00394779423238312,-0.00422457465385673,0.0120247781192235,0.00508608309389769
"1639",0.00719724914002473,0.00279613500057274,0.00520814531012448,0.0131050461310511,0.0010253278602268,0.00168093302058447,0.0127043362267061,0.00798625030288513,0.00928793390866134,0.0062280993616175
"1640",0.000363130431931147,0.00709748371972152,-0.00345430650098744,-0.00950356185586343,-0.00782138254972453,-0.00355471447952693,0,-0.00594201202172995,0.00273581488801655,0.00309481492883301
"1641",0.0136211762943714,0.0279388806029683,0.0294628173394231,0.0490404592729916,0.011730689235365,0.0100083231955281,0.0276283634189962,0.0328763121744742,0.0272013318032576,0.00501346891729848
"1642",0.000417413573514658,-0.00759085164296125,-0.00168334029271122,-0.010670785508596,-0.000834898390411509,-0.000785269726336191,-0.00653941561449167,-0.007957406035354,-0.000885391192617324,0.00383732509349644
"1643",0.00382096204745186,0.00444140859541808,0.00927470612024051,0.0102722758892468,0.0052916807109129,0.00314220296912948,0.00365671772927723,0.00607686714958389,0.000402827690393126,-0.00267588302880972
"1644",-0.00374665444860911,0.00122806480081739,-0.00835413462407975,0.00406716685150488,0.0034162634679078,0.000489540217296414,-0.00160336921838855,-0.002657823435536,0.00571749879207606,0.00114992905154732
"1645",0.00256711715495483,0.00147204673455659,0.00926696323329801,0.00911411544478091,0.00184077930302151,0.00440165210845223,0.00525575396278666,-0.0031489972435963,-0.0125710546286417,-0.000765765091293669
"1646",0.00547750150946325,0.00857422935580243,0.00500825983278563,-0.0117915333187582,-0.0124926394066947,-0.00467508310256082,0.00624459421561752,0.0026730832157269,0.00559521569899446,0.00421458075059888
"1647",0.00177669337149333,0.0029147740549107,-0.00747507963978211,-0.0027923130298636,0.0158133968151386,0.00548057113474232,-0.0010105133674736,0.000969545160759422,0.00887024419207738,0.000763017835870849
"1648",0.0019507242143062,0.00484389615122538,0.00251054399534723,0.00992845592417546,0.00146541960449986,-0.0000977751521776815,0.00288933892731125,0.00508482105265973,0.0298137236846479,-0.000762436083540319
"1649",-0.00212406677543031,0.00168705522918611,-0.000834713821576627,0.0108393586651712,-0.00420648088869424,-0.00116786313178996,-0.000432080800389478,0.000481545259870986,0.00675264690321775,0.00152611420787818
"1650",-0.00366531124884484,0.00288750819650851,-0.00835413462407975,-0.0102242656853181,-0.0126718536446839,-0.00672364285863214,-0.0194551023874096,-0.0086683916466419,-0.0171922278903276,-0.00799996926074609
"1651",0.00243272057103128,0.00575804373938116,-0.0185342761272566,0.0057947986057485,-0.000372145519264899,0.00147156349392286,-0.00117595680108629,0.00364344971368058,0.0093347581737977,-0.00115205797759044
"1652",0.00106561699061292,-0.00238549227979767,-0.0231759545339051,-0.0022543614143179,0.00614071482218637,0.000881604934367175,0.00264882374614328,-0.000968171686319574,0.000854907917228864,-0.00615151468866593
"1653",-0.00307501211335826,-0.00382604624272109,-0.0219683520503358,-0.0125533745161952,-0.00730509258425183,-0.00205580979619668,-0.00792493008842865,-0.00823628313285363,-0.00240719057623229,-0.000386841912370151
"1654",0,-0.00336054411194509,0.00898461093266034,-0.00228817941574921,-0.000373500225038681,-0.000293729333673665,-0.00118361100719955,-0.00610655365850821,-0.00272441813089119,-0.0034830042132139
"1655",0.000711979676581542,0.00602143102746378,-0.000890460650768143,-0.00586139877329483,0.00363483400529274,0.000686540059984919,-0.0137735783288175,-0.00442365288958046,-0.00124879805060862,0.00699035586535879
"1656",0.0115581783899779,0.0100547645666818,0.0276294004909297,0.018200080418912,-0.0192684427729715,-0.00882604194366043,-0.00555646472254623,0.0118488928347293,-0.0105501563812922,0.00231393010372782
"1657",0.00169897245283646,0.00568875389511692,0.0156116315553585,-0.000251642604873759,0.011009981917292,0.00851833539242963,-0.00437905936754102,0.00146393199978401,-0.00197456755410652,-0.00384769978730604
"1658",-0.00146237722033871,-0.00259270169804648,0.0025617140745906,-0.00629543792781184,-0.00769793802045393,-0.00314263317428487,-0.000606981304382082,0.000487079669117652,-0.00522320350408989,-0.00502117525665891
"1659",-0.00568207986909219,-0.00165396836227627,0.000851801383985773,-0.0126711986506385,0.00293276059448999,0.000295505759437598,-0.0034905720067282,-0.00146108037310133,-0.0137628961120818,-0.00815226196392715
"1660",-0.00324078735667788,0.00142044539343256,-0.0187233990044424,-0.010780370830044,0.00745251761830135,0.00364372257430845,-0.00411219772244642,-0.00658361718678746,0.00145197223963889,-0.00665361032499945
"1661",0.00366485717270981,0.0103992262106134,-0.00520379719143449,0.0192011272250223,0.00271451684081647,0.00147218823325446,0.000917616925767639,0.011291074119663,0.0218284249403395,0.0051221547324638
"1662",-0.00288548726559956,0.00163710718691479,0.000871828350458959,0.0020363954578464,0.00158778264360193,0.00068614746905582,0.00947276507011496,-0.00169891682515522,0,0.00705608126312685
"1663",-0.00118141970448593,-0.00373647143275058,-0.000871068927872365,0.00940059558308892,-0.00680589284401134,-0.00195828644111495,-0.00817314569911776,-0.0070504363651529,0.0178937725217267,0.0120669074580908
"1664",0.00295647482936645,0.00609471032317899,0.00871828350458803,0.006040572233313,-0.0144560805363559,-0.00902693091504547,-0.0137339053770204,0.00171368328821808,-0.0107643998000311,-0.000384530976713426
"1665",-0.00512949623609193,0.000233217588825108,-0.00518573526885902,0.00325239323154891,0.00152399224532029,0.000890838518383008,-0.00216642960448465,-0.000977597117130857,0.00986380162617517,0.00807999927135161
"1666",-0.0139856775067201,-0.0051247301667271,-0.0139009451850375,-0.011471361044767,-0.0135044897985468,-0.00553969622454131,-0.018917487953954,-0.00905336667690337,0.0208527286821705,0.0095419721382568
"1667",-0.00330562035176563,0.00210711640196637,0,-0.00857695749435483,-0.00347083716806407,-0.00387904073497192,-0.0230758973104827,-0.000740506560158671,0.00675829589553811,0.000378066669932675
"1668",-0.00639234834161162,-0.00887840207759238,-0.00264325967685353,-0.0188296871468735,-0.00870632631856993,-0.00429387299310058,-0.0135900412408417,-0.0113667865507208,-0.00429934372757068,-0.00113377136863213
"1669",0.00491603219109216,0.00353596343087847,-0.00883400487638997,-0.00181520731708229,0.00770961917504143,0.00541563296433822,0.0234542931748214,0.00324934294666313,0.00333309610382138,-0.00189184165773648
"1670",-0.00616028645440758,-0.0112755804436938,-0.0142600684421138,-0.0233826622253877,-0.0109431213945713,-0.00628430591626006,-0.00208334695979095,-0.0174390464050673,-0.00286893173731062,-0.0011372096858524
"1671",0.00911498054440774,0.0125921977248018,0.00632903237831184,0.0162275796108744,0.010183029055659,-0.000401710252976417,0.00562059690032379,0.000506891129139042,0.00560302082818853,0.000379579586898826
"1672",0.00337240419440832,0.00610042974417291,0.0170709596566356,0.0117801489108056,0.0108557896877199,0.00562377763026634,0.0116575919906952,0.00734943378131225,0.0157367369284953,0.00796658499444414
"1673",-0.00372084959008978,-0.00629665154143932,-0.0114840010155703,-0.0108665981739087,0.0049862390272688,0.0019972566141786,-0.00378821743938051,-0.00654087124497804,0.00407711656384513,0.00564542635091381
"1674",-0.016084160805488,-0.0194789174906257,-0.0107238460716564,-0.02301866295041,0.0125940245620235,0.00568081368670281,-0.00301083967975924,-0.0157002682079449,0.00959765986558136,0.00973052179638567
"1675",0.00355075402795979,-0.00215436397626045,0.00271021710531438,0.00214174673761436,-0.00810307333221993,-0.00406311374075996,-0.00476797046182442,0.000772143579793827,-0.000292453382084168,0.00148263579272623
"1676",0.00158639149170647,-0.00263829147557737,-0.000901188243820683,0.00801518693605385,0.00797943661524592,0.000994835603807642,0.00159696505294549,-0.00128573068366544,-0.00614448070359619,-0.0103626668671772
"1677",-0.00316754177556444,-0.0108227670803879,-0.0198378618561539,0.00768583624855457,-0.00113107792198397,-0.00188830682463281,-0.00765276283749283,0.000514844801336567,-0.0091999708986521,-0.00299180861046588
"1678",0.00452206542140976,0.0143450293797505,0.0248391764768532,0.00631274278204219,-0.0141037475978312,-0.00567555837743949,-0.00835491192733495,0.012863474735906,0.0133709929197368,0.00525124106240105
"1679",0.00827281563695981,0.00479385597242055,0.0152602273073033,0.0177729676250142,-0.00220700275055452,-0.00331023199461855,0.00712893219925381,0.00457211356342269,-0.0129012903225523,-0.00858201128343494
"1680",0.00126711309053684,0.000476875322934944,-0.00265251067899708,0.011813086161315,-0.0139441853655841,-0.00764928428520517,-0.00852637684204494,-0.00176993779172352,-0.0182682825406718,-0.00225815504595728
"1681",0.00048210149956196,0.00643800790749616,0.00354617688207148,0.0147209256615468,0.00497355020894141,0.0060858048469814,0.0183351783488284,0.00329278359926244,0.0147503558566646,0.00565820345158907
"1682",0.00957592440058019,0.0106607785461648,0.0256183648198507,0.0262630738404408,0.000484881007786431,0.00201604004708034,0.0197578547609021,0.0217119050409662,-0.00178896765362513,-0.00637662282010609
"1683",0.00739707128298872,0.0128927753822412,0.00775193428949672,0.00755533972736067,-0.00698270619852082,-0.00462795424198048,-0.00125004835694331,0.0113663658352079,-0.0162049057962839,-0.00906001565387571
"1684",0.00313847851672655,0.00740549267210411,-0.00683751951668155,0.000725762885528836,0.00888841422644804,0.00505359917642245,0.00688373013768451,0.0046420363851567,-0.000303689073034463,0.00152390635694055
"1685",-0.00265613846143276,-0.00413509556470015,-0.00688475974170399,-0.011602529548285,-0.00135544068161408,0.000100749827011803,-0.00637047732028806,-0.00583669677874921,-0.0305998412437321,0.004944778001164
"1686",0.00224891349425183,0.00392180392689956,0.00519938417631205,0.00660298716115459,0.00387758300465491,0.00130706442222839,0.00218908358169601,0.00660479524461399,0.00117491973329531,-0.00302796768043412
"1687",0.00578749961637848,0.00597416143765428,0.0129310352024701,0.011175936633522,-0.00666350923080905,0.00220902647186794,0.00983009207974539,0.0080192496471807,-0.0107182209356907,-0.0125284973465647
"1688",0.00446283091026256,0.00137050318536391,-0.00425540572827832,-0.00216239116001926,0.00826370823040934,0.00200444488949136,-0.000772523907001887,0.00699152872112618,0.000395436940975102,-0.0103806785639978
"1689",0.0115738401899543,0.0253193894937807,0.0307693108134122,0.0418974376241923,0.0123419081989526,0.0123996552431906,0.0349465378145997,0.0277710293738997,0.0435572727272728,0.0217560449952168
"1690",-0.00167591122300226,-0.00489435140566452,-0.00497522106026338,-0.00531549188905167,-0.00590514957592669,-0.00345718808056661,-0.00388475788947529,0,-0.00196950996021172,-0.00380226857225308
"1691",-0.00699149916626673,-0.00558920215377201,-0.00833331930627246,-0.0223048100919977,0.00526999094572211,0.000991563718008903,-0.017249020059887,-0.0112541678078772,-0.0287666110056927,-0.0091603372497493
"1692",-0.00462730674098633,-0.00382184803626051,0.00336141788891897,0.00356447828393947,0.007338762699582,0.0037623979857444,-0.0064103570565559,0.000237029559334134,-0.00320409505473651,-0.00731889206234926
"1693",-0.00235393483703694,0,0.000837440663423061,-0.00852440668909249,0.0107861100802857,0.00365031682193084,-0.00660496970541757,-0.00189682310285688,0.000862414719033699,-0.000388042802127453
"1694",-0.00289040027079435,0.00225685053868618,-0.0025104513767078,-0.00764278614387581,0.00205967247856176,0.00275206568767317,0.00343368266098754,-0.00237524187690041,0.00885155071748245,0.00155269384311052
"1695",0.00384535205823888,0.000675611598614623,0.0159396723679954,0.00409150841296846,-0.00700630190219353,-0.00215628247118582,0.00606634664872008,0.00499995099929884,-0.00776451630057939,0.00775195220958547
"1696",-0.00459676781909035,-0.000675155455757914,-0.00743177905128478,-0.0117450184593179,0.00244613147052486,0.00137513784266963,-0.00371056577253537,0.000237005379424282,0.00923389929388918,-0.00499997149863052
"1697",-0.00532826481836535,-0.00653018304267816,-0.00831963616174847,-0.0113994986477234,-0.00150148794600302,0.00166779621470381,-0.0100868901841568,-0.0021316081480216,-0.00612551751472812,-0.00425197135461264
"1698",0.00791642213031274,0.00770617406369589,-0.00419446125447809,0.0198724506823325,-0.00303450486868984,-0.00222621017912139,0.0152062130927848,0.00688346250567129,-0.0280074675928559,-0.00659936835062425
"1699",-0.00094509761295114,-0.00134932626337358,-0.00505483436749365,0.00384876326547712,0.00151232124211242,0.00167027543948639,0.000617611086776826,-0.00117869499247536,0.0198250427747024,0.00976938764059976
"1700",-0.00922094204884161,-0.00495487170171172,-0.00762065615230845,-0.00383400707986847,-0.00160457244990941,0.00137386017369523,-0.015432262682139,-0.00873272255820257,0.000944451455130668,-0.00154804612847681
"1701",0.00757707551716114,0,0.00170646268440877,0.0129898396957406,-0.000755885954198621,-0.00274386147034644,-0.00360488042581686,0.0030953675811094,-0.00511087435131308,0.00310081279751295
"1702",-0.0086450464151776,-0.00520597524735833,-0.0187391590709212,-0.00854869887457277,0.00406760361591552,0.00088468114953244,0.00440470930698389,-0.0113932745622617,0.00877262316266991,0.0069552021763386
"1703",-0.011646463219254,-0.0102390412972611,-0.00347239310692171,-0.00958103200403826,0.000282500200811775,-0.000491047663760513,-0.0114331824555356,-0.00384144677528009,-0.00188026482200143,0.00345352149477884
"1704",0.000725307432946076,-0.00275862209656097,0.023519150284071,0.00749698216060835,-0.00800579242884003,-0.00176789679810241,-0.000317132169727175,0.00964095675782772,-0.0101255963873533,-0.00726575415014186
"1705",0.0215577769656854,0.0205164166441045,0.0144679932761642,0.0235238173180525,0.00161397501394966,-0.00216528269006344,0.023930485572337,0.0181424284291265,-0.0145904685227938,0.0127119685621264
"1706",0.00644316424945313,0.00609894792735144,0.00167792377940001,0.00445584640259944,-0.000284408929857927,0.00147910949433738,0.00959628415028702,0.00281343453743488,-0.0134384730048719,-0.00532534128258155
"1707",0.00399390701725522,0.00291862061211412,0.00167513624140159,0.00583716276224044,-0.00805969020412067,-0.00334818660338021,-0.000306815150598605,0.00327334577867622,0.00187605223288823,-0.000382403970200285
"1708",-0.00725379808421178,-0.00268636818548884,-0.0083611190163132,-0.00974937818661881,-0.000669278505797011,0.000197836327931356,-0.00322039611723146,-0.00838952471328447,0.00732720821741917,-0.00344303107689314
"1709",0.0139656620429149,0.00718293555562655,0.00927470612024051,0.00796977352892436,0.0125311807249637,0.00484086865381772,0.0181537886584859,0.00846050432339251,-0.00153561784040357,0.00767759687630321
"1710",0.00668318622665298,0.0147093952544932,0.00835401904423039,0.00627930363834484,0.00906923787077063,0.00570145930606003,0.0154125130452076,0.0139829572935,0.0314068072575133,-0.00533326056285455
"1711",0.00675438188536948,0.00636925546674316,0.000828604552449042,0.000924414822592423,0.00215327064390713,0.0000976198536080108,-0.00193448754681935,0.00873368019458365,-0.00447339514163236,0.005744925346165
"1712",0.0000573454583125965,0.0015277070154629,0.000827804007986988,-0.00161593882907751,-0.00317616999945636,-0.000684138441023552,-0.00521839047931827,-0.00273397992497049,0.00102487191209888,-0.00228489091290041
"1713",0.00579150045114307,0.0126390519271182,0.00496287609754931,0.0097127667800867,0.0111526469469703,0.00694443418099722,0.010641626256527,0.00525435968316423,0.0185855484662416,-0.00114502251469084
"1714",-0.00478883808990649,-0.00602550684524195,-0.0205762090047192,-0.0233622006975779,0.00389308632996199,0.00174806072702549,0.0020761019851121,-0.00659075685163879,-0.00502546791481284,-0.0152846645628761
"1715",0.00332252834297542,0.0073609259099976,0.0100842071628604,-0.00211074526170762,-0.00387798898406044,-0.00203582153125148,-0.000739776457556296,0.00205891302072869,0.00940237766100904,0.000388042802127453
"1716",0.00456746283691833,-0.000859772519551827,-0.014975032021709,0.00470036708814048,0.00370774924872053,0.00174933180260806,0.00977462865673662,-0.000228047756405503,0.00431110874416207,0.00310321811263736
"1717",0.00159115184855096,-0.00408691783636539,0.00337828789945305,0.00584776208281812,-0.00341732494881941,-0.000970199183237819,-0.00689351290996987,-0.00411068884361299,0.000766449445307904,0.00386688312838346
"1718",0.00533403038374036,0.000648058630437598,0.0075757533410139,0.00325609025050366,0.00129775483038208,0.00135908833712395,-0.00841823386202967,0.00114627311903726,-0.00605081197994506,-0.00269645895743109
"1719",-0.00496676020454168,-0.00366934131024177,0,-0.00556330971407748,-0.00601497300230069,-0.00261734318973939,-0.0072981713477811,-0.00847412317185003,-0.0013099945654621,0.00308999375752017
"1720",-0.00283678257141473,-0.00498256539859021,-0.00501262871665498,-0.0102564520467331,0.00214157149084548,-0.00116668074991788,-0.00720172530143481,-0.00323405766195872,-0.0143519129158065,-0.00847131645656707
"1721",0.00238983972376849,-0.00631396941287843,-0.0109151045590405,0.000471024852145119,-0.0108250194308196,-0.00554679399778424,0.00634703985561047,-0.00324464872903574,-0.00618444506316651,-0.0124271349969011
"1722",0.00351832661497298,0.00591587228183776,0.000849002971733404,0.00612073896584109,0.000941632031749906,0.0019609257625246,0.00135183852107668,0.00278975457625652,-0.00110278852546963,-0.00432562145749138
"1723",-0.00316705892203262,-0.00936627465644813,-0.0084818655471447,-0.0201217802099829,-0.0119480210756774,-0.00450064447822718,-0.0151471930232391,-0.00765104589568621,-0.00197145338650662,-0.00276465649222335
"1724",0.00510588452990346,0.00945483120231949,0.0136868306564424,0.00310395230403859,0.000476178912561576,0.00304620262367372,-0.000151913598553266,0,0.00505688219116451,0.000792149946476695
"1725",-0.0126434184192837,-0.015465070467779,-0.0185654906184489,-0.0180906468869231,0.00847066957850662,0.00264572738260194,-0.0121842493629626,-0.0135513182086211,-0.0081760457903155,-0.00712309554301804
"1726",0.0134913492775723,0.00553097805901825,0.00773879441853786,-0.00218209430706484,-0.0240658314359892,-0.0112371072989794,-0.0134132176394359,0.0045002656789388,-0.0149017512713459,0.00557991813609582
"1727",0.000169324979420127,0.00308031374899875,-0.00170658072969698,-0.00510185632187232,-0.00377167780235965,-0.000494081447939387,-0.000781542714727079,-0.000235621762755933,-0.00329897009413405,0.00435987023310913
"1728",-0.0020302403013035,-0.00592257090591186,0.0128205146396987,-0.00537255357740329,0.00465941965670402,-0.000889730155375412,-0.00344082326800721,-0.00165090464640993,-0.0114636793865259,-0.00670879114630474
"1729",0.00802435414018432,0.0044132948327138,0.00759500315307493,0.00171883709425935,0.00367145452730244,0.00415639272052615,0.00706216954039296,0.0011810676982531,0.00326664769130214,0.00437042702655299
"1730",0.0049896228421209,0.0024165190128973,0.00837512502979609,0.0161763221232361,0.00616108119535075,0.00482875901577451,0.00794767896947546,0.00802263090978483,0.0115588036069809,0.0043511245202319
"1731",0.0043509233470993,0.00416383917135721,0.0141195821076014,0.0190546557783398,0.00200908129913713,-0.000784371158518038,0.00247363820429691,0.012406110206348,0.000402373873075623,-0.00157540193747197
"1732",-0.00349921806321518,0.00240080209590987,-0.00163807142312289,0.00899392584692538,0.00601509143778212,0.00353325931389037,-0.0069402417818214,-0.00346806276552192,-0.0114221203346203,-0.00670606351599057
"1733",-0.00217379249477878,-0.00239505204992851,-0.00574224828486836,-0.00609898552417576,-0.00759269172242338,-0.00371695482483347,-0.00760972725430231,-0.00719217921358917,0.000406794134958588,-0.00158862234773016
"1734",-0.00312793766903063,-0.0104758061977032,0,-0.0136888444427538,-0.0170238071045685,-0.00549693650854921,-0.00876368453626142,-0.0100494980488829,-0.0230174385445491,0.000795534102772777
"1735",0.00806872921921875,0.00992514195437089,0.00412549658987782,-0.000957125435392392,0.00165442431429863,0.000887988523022631,0.00536776862616417,-0.00165249725449002,-0.00149850978608446,0.012718632235597
"1736",0.00500238329044067,0.00502293061648729,-0.000821773019853089,0.0071853871050096,0.00932448525277874,0.00286047825868274,-0.00298340734680458,0.00118231846748396,-0.000166783388914737,0.00313971495238485
"1737",-0.000995573576284214,-0.00173867933385607,-0.00740149386062294,-0.0128416456783353,0.00288756043736083,0.00078627427504685,-0.00425276736865443,-0.00661291152748045,0.00450301041532697,-0.00117365263192004
"1738",0.00027682836359233,0.00152382121820271,-0.00414222040619749,0.00337263281551858,0.00374238368235003,0.00216188198716516,-0.00284733417402261,-0.000713451113986463,-0.00531295870258142,-0.000391771302957644
"1739",0.00243508289737027,0.0036949663322956,0.00415944976388816,0.00648238938648338,-0.00172131412862364,-0.00225506894697336,0.010310983026192,0.00499638190259066,-0.00300451510599231,0
"1740",-0.000662481427646244,0.00346471371518486,-0.00082830653448851,0.0102575713250397,0.000287513912400339,-0.000589768417623482,-0.0092638912104277,0.000473373736791238,0.0103800268741003,-0.000391844188296631
"1741",-0.00259663232462659,-0.00798428756757363,-0.00248757611493755,-0.0210151345879274,-0.00777798612235558,-0.00429440173673745,-0.0052297014536975,-0.0134880870496825,-0.0258491721420673,-0.00117599337105756
"1742",-0.00432065882847799,-0.0100066291041776,-0.0041562686348624,-0.00337670046623118,0.00367751971812846,0.00178072946689567,-0.00111504434633636,-0.00407765667367643,0.00323181658051008,0.00588701097795474
"1743",-0.000111175975896383,-0.00549340805262788,-0.00751260916758756,-0.00121024589224372,-0.00954583664329278,-0.00454279678130409,0.00223286293060387,-0.00192660212203266,0.0169549001098246,0.00195089246041613
"1744",-0.00439533581543172,-0.00397693100750562,-0.00841022858947127,-0.0058152799830804,-0.00282305112785286,-0.00247966440061176,0.00111396447919065,-0.00506734795966202,-0.0138379127529001,-0.00116836855358804
"1745",0.0111768609386094,0.0135314278478669,0.0127225284285621,0.0221788872351829,0.00478358506727927,0.000894545053452545,0.00778887184220522,0.00654851046250871,0.00211327129044969,0.00350880445250534
"1746",0.00254232398566856,-0.000437737140972727,0,0.00143067734821378,0.00233181080880795,0.00119282344933591,0.0064668744678078,-0.000963934862336813,0.00986923635927694,-0.00349653579214948
"1747",-0.00358315359303885,-0.00394112322734064,0.00167513624140159,0.00047618367382829,0.00717352976787167,0.00416808745785358,0,-0.00241197532728288,0.0175409203346064,0.00311894620786823
"1748",-0.0112311088185472,-0.00681480751162811,-0.00919748309266799,-0.022132386347068,-0.00769999550808997,-0.00385440178591057,-0.0216265911332877,-0.0159574172591587,-0.0078804711869972,0
"1749",-0.00330143494367263,-0.0108456199937736,0.00337550766235628,-0.00584075419881425,-0.00378241394451839,-0.00287704171985192,-0.00672759924700417,-0.00491409851976832,-0.0212642725362876,-0.00932762588406888
"1750",-0.000111989046382877,-0.000447532130515294,-0.00841022858947127,0.00244805840814188,0.00486821895063705,0.00149270552106673,0.00403160454433871,0.00197536733809889,0.0092146080884723,-0.00392313431467806
"1751",0.00623166314956003,0.0123126438929264,-0.00593732231121935,0.00659339637593104,-0.00368230679749171,-0.000496995653735066,0.00112440334065922,0.000246351620043272,0.00259679182267036,0.00315080387494393
"1752",-0.00318004137377415,-0.00457720944830442,0.000853042469743492,-0.00873391890871733,0.00447397747464207,0.00318055726919497,0.00529438704601248,-0.00812989326142133,-0.00868911339812661,-0.00471136123717364
"1753",0.0170723451721642,0.0156250678515926,0.0195843596584198,0.0199042973570234,-0.00503458737054385,-0.00376519663922226,0.0175549052125341,0.0116740910980002,-0.00876528430231294,0.00197235968110299
"1754",-0.00115581223071648,0.00307697820290587,-0.00842440523321475,-0.0184020221298921,-0.000973132514868857,-0.00417643141954038,-0.012233385473437,-0.000491200152554883,-0.0237224808798361,0.0023622536040393
"1755",0.0058168447915643,0.00328649997859531,0.00339834018932472,-0.00147985747201518,0.0153889234167062,0.00309545701909375,0.00778031665841006,0.00326208048367294,0.00975441560703727,0.00785547348507354
"1756",0.00534256274167277,0.010919357534348,0.00931406896759879,0.00741104440324669,-0.00565930185251518,-0.00318586214939875,0.0014155172882262,0.00825448483206914,-0.0031913230431031,0
"1757",0.00219153298963337,0.00691319724930439,-0.0134228359550707,0.00588526475980555,-0.00800719780212,-0.00389498493414753,0.0017467767012902,-0.00173654695557102,0.00458594791035738,0.00311765026524369
"1758",0.00508391997037649,0.00493435835365585,0.016156482065093,-0.00853253166551993,-0.003853626457892,-0.000864220269060856,0.00110980531638361,0.00372777264170199,0.00551248932838044,0.00155406033549488
"1759",-0.0000543750655374042,0.00533736705027787,0.00502103894533423,0.0154905634686311,-0.00284004907263047,-0.000602649692397428,0.0012666855828356,0,0.00325513968228774,0.00271524598323292
"1760",-0.000163060200582765,0.00339772294065455,0.00915905475772538,0.00435820754362815,0.00687522266445462,0.00271548088628504,0.000790691939788868,0.00940819844311069,-0.0147712086380325,-0.00580270831542484
"1761",0.00473286001511264,0.00423289818828421,0.00164997712953463,0.00771484612167206,-0.00634102580033025,-0.00451383235387537,-0.00316044869316878,0.0105465856579214,0.00632640615587476,-0.00155639897877735
"1762",-0.00958363352412261,-0.0229716857382819,-0.0164743563555104,-0.0385167687538027,0.00304323957549113,0.00392966844017129,-0.00158530451641903,-0.0189319910207802,0.0161901218690117,-0.0144193330254777
"1763",-0.000164167624208011,0.000862960684752112,0.00586270400886524,-0.00174172042647325,0,-0.00060209405486511,0.00587497238488099,0.00544268725885799,0.0109322118644068,-0.00632664688813733
"1764",-0.00289800493839887,0.00172422747178036,-0.00333068177587947,-0.00947162789594769,0.00420889160031335,0.00281197601205685,0.00410396089178411,-0.00344465593487686,0.00176040739575489,0.00119377599891823
"1765",0.00614182060371826,0.00709963104823497,0.00417735713167433,0.00427763815860294,0.0025342838614808,0.00160212578936858,0.00345848394815973,0.00172860496601634,-0.0056903765690377,-0.000794901731337117
"1766",0.000218351644983628,-0.00170909997124435,0.00166386382097339,-0.0032570721602414,-0.00272195300184808,-0.00489917140558638,-0.00156653903506421,-0.00419027165733554,-0.00589123884867859,-0.00954649111203931
"1767",0.000653579947207383,0.000856025767816071,-0.00332238242692806,-0.00527915881610541,0.00584899104136727,0.00261263951062141,-0.000470788311053183,0.00173281499048383,0.00287839477958696,-0.00803205995609246
"1768",0.00272264505204367,0.00962159382112371,0.00666675469838185,0.0176900769625659,0.0119207534938413,0.00841868305145543,0.0119310247809576,0.00716567581040684,0.015195027985776,0.00647764372042814
"1769",-0.01330505196133,-0.0084711242005906,-0.00662260342587684,-0.011919513575515,0.00498019626472423,0.00288165053704459,-0.00651568777419853,-0.00662417040032359,0.00631959909663071,-0.000402247119002164
"1770",0.0108977829328305,0.0128149909229103,-0.00250009308552912,0.010806914832306,-0.0045741970067088,-0.00376556554206187,0.00624623869897811,0.00419844853013918,-0.00933728332516814,0
"1771",0.00538996284542415,0.00421774917933382,0.0075189170527592,-0.000248676275743098,-0.00105307814108246,-0.000895050015314314,0.00465540293271416,0.000245763339677518,-0.00191838353422624,0.00281690432515114
"1772",-0.00129975249410952,-0.000209956610136786,-0.00331662251152542,-0.00547121515160165,0.00670860559113096,0.00278752865530985,0.00231690553211705,-0.00122912546949305,0.00108638639189751,-0.00160515579427789
"1773",-0.00422934031056532,-0.00483101887592197,0.00249568149589741,-0.00500144410994274,0.00418880920984543,0.0023829074656927,-0.00323609973562489,0.00221547464540084,0.00951664571736677,0.00120581268813291
"1774",0.00294061540419333,0.00548753134695801,0.00165972168427775,-0.00150775113746604,0.00075885174832635,-0.00108963910534199,0.00695710512964065,0.00343920660277242,-0.0101711982138428,0.00240863827526017
"1775",0.00065152681081293,0.00125941132504148,0.00248561662625102,0.0133400330561615,-0.00246356318312968,-0.00277627525846402,0.00261035792461528,0.00416127964001856,-0.00426060996476041,0.00480578379051
"1776",-0.00819302774572472,-0.00167703621381354,-0.0198348121820553,-0.0245903452859302,0.0141503163541179,0.00676138004837457,-0.000459488492525639,-0.0107264226701915,0.0218139018069652,-0.00079720148395801
"1777",-0.0213359289622417,-0.0317092879170057,-0.0151770523348445,-0.0262283736580906,0.00646147623958293,0.00404923402241009,-0.014708183807011,-0.0197140417008947,0.00410542734128061,0.000398959814302602
"1778",-0.00491956950583161,-0.00542202168270289,-0.0128424502933567,-0.00392274582579388,-0.00697857702578497,-0.00304894026306357,-0.00606418590669144,-0.00351922840454166,-0.01087580332917,-0.00677829885603132
"1779",0.00595480761928213,0.010902874259501,0.00867311158203132,0.00630089483621843,0.00243672303947262,0.00147976197032929,0.0101685487789813,0.00983825728883336,-0.0000826884927470628,0.00481735918529047
"1780",-0.00960514311482297,-0.0138048994695855,-0.000859900778935718,-0.0143490338441313,0.00822485876717982,0.00472893450401823,-0.00464587523934101,-0.010242291902958,0.0125672099024525,-0.000799030209567286
"1781",0.0106007050677617,0.00393679481998976,0.00172097445265562,0.00926427781398931,-0.00287385761187742,-0.000980709679201941,0.0121364310795513,0.00706719503316444,-0.0220462478807361,-0.00399842815131779
"1782",-0.00585877639585786,-0.0137254264130815,-0.0266321894469745,0.00157339101224196,0.00669385686013957,0.00392632342994226,0.00307435572905979,-0.0105264177160646,0.00267177931047291,-0.00120436045501515
"1783",-0.0225051039845126,-0.0203225140704832,-0.020300166346488,-0.0282796919684274,0.0121845676485308,0.00543597438739596,-0.0145591678764526,-0.0167170344725773,0.0102423519108119,0
"1784",0.00700428409516429,0.00901909764458209,0.000901132483273948,0.0202103240044194,-0.0106109242741762,-0.00301970288210873,0.0104198851418438,0.0118495560566281,-0.00272009561490272,0.00763659306640951
"1785",-0.00125404099484416,0.00402244963123244,0.00180004910573128,-0.00369794103753229,-0.00924569859075075,-0.00361519642778629,-0.000308004748738711,-0.00152729864540857,0.00247956860037313,0.00199447064194791
"1786",0.0131870808952297,0.0213667269439997,0.0116802334956105,0.0209436636374025,-0.00429267928100152,-0.00186338723440838,0.00739028607640591,0.0137678395098582,-0.00041225986963267,0.00398087837775551
"1787",0.0123959584177427,0.012421079702134,0.0159858724133979,0.00571297687765493,0.000843732312646228,0.00265246477410241,0.00672485514829702,0.012575832173612,0.00767073585732003,0.0114988169728101
"1788",0.0018363914506474,-0.00258310370370662,-0.00437079147033703,-0.0111025689398977,0.00280904911341073,0.0004901385915832,0.00910896194251043,-0.00571306951233119,0.00613898675843472,-0.00548796906493509
"1789",0.0109440408775989,0.015105909111057,0.014047402853854,0.0216711016917601,-0.0057891244645889,-0.0044069970709224,0.00345992657777505,0.0174870441317148,0.0117149611408225,0.00512409213369813
"1790",0.000494574220003763,0.00276359674195947,-0.00173157114081068,0.000255515701197195,-0.00516612846428177,-0.00236089797194439,0.000599956400566315,-0.00147333306118391,0.00056287390991594,0.00196075756439518
"1791",0.0051625629965999,0.00678394572701713,-0.00867301630975614,0.00102191857587663,0.00566458664838088,0.0047330590361323,0.00389544697350819,-0.000491609474797206,0.00851882986418051,0.00547949829681849
"1792",0.00551914614093829,0.00547461871072863,-0.00437444781209861,0.0122512335066107,0.000563431390164792,-0.000687397451970551,0.00402997893447088,0.00368990287719417,0.0132281777548517,0.00350334094595328
"1793",0.00119541411052215,0.00607356540452497,0.021968434938447,-0.00932949930542448,0.00225197418759238,0.00245530832734508,0.00594611587157057,0.0095587481817847,0.00196618164425977,0.0143521342519306
"1794",-0.00662164179809943,-0.00666126285837132,-0.012037973346854,-0.00687193694439225,-0.00421306800746313,-0.00195907517967175,-0.000295435445795689,-0.0024276190610506,-0.00886974083406999,0.00267682779140133
"1795",0.00590077584642579,0.00586756618006889,-0.00609221837615492,0.00358800816403715,-0.0024438443552095,-0.00107981299977822,-0.00177393977616147,0.00803119567166166,0.0105329930434701,0.00190703312623652
"1796",-0.00114059066733163,0.00166685290582569,0.0078807713886615,0.00689463201147733,0.00527764129744157,0.00127754329452578,0.00162897470070233,-0.00193129733050956,-0.000156708466406141,-0.00266463921158044
"1797",0.00554691465034796,0.00665542287086551,0.0112945193056191,0,-0.002531381876687,-0.000981572280831067,0.00162645623929381,0.0024188097605522,0.0110519123522197,0.00419845517025497
"1798",-0.000378690478715749,-0.000826390644169006,-0.00343629509873367,-0.0114124369315098,0.00892887835565248,0.00343796930940976,0.000442573805715218,-0.0024129732373338,0.00170557400939697,-0.00456098027062002
"1799",0.0000541847331678724,-0.0047560958093017,-0.00431033972535777,0.000769643570279976,0.00530958896381861,0.00293673759080915,0.0028030325799191,-0.00362878206046091,-0.00851331894131058,-0.00267273931650935
"1800",0.00524738156668758,0.00540201989152056,0,0.0189692573666882,0.00546668920048998,0.00117163876640292,-0.00102968339122844,0.00194265133533955,0.000702490042131743,-0.00306282394495516
"1801",0.00252918932156554,0.00289321179485857,0.00519473719925823,-0.00679252792586793,0.000553184506777216,-0.000975072636903218,0.00662712544106814,0.00508808884626544,-0.00452413427123555,0.00345609488391885
"1802",-0.0070322783406207,-0.024727177680151,-0.0232556412246436,-0.0177302915576182,0.00667517274606877,0.00494624519117348,0.000731813845386897,-0.0106070379916682,0.0209214068111252,0.013777356550581
"1803",0.014056150833244,0.020283371371127,0.0255731977922884,0.0170188944125849,-0.0150418875058651,-0.00768427970091956,0.0122807928353497,0.0160815167943791,-0.0123570503223529,-0.00377495795619198
"1804",0.000906038077092219,0.0012422612932097,-0.0111780017281133,0.000760899137216553,0.00214173108517168,0.00107835188650274,-0.00129986163463869,-0.00311739272920952,0.00163200195387003,-0.00833649397690217
"1805",0.0022903652178794,0.00868671854690772,0.0191303814570809,0.0141880258238427,-0.0098495435658057,-0.00430875015141186,-0.00477227136267833,0.00793832696299712,0.00993094118962645,0.00917079873772564
"1806",0.000425050383246584,-0.00676636732518721,-0.00682612226336032,-0.0127404587740887,-0.00628699583377523,-0.00432629874096579,-0.0113338161021139,-0.00119324110616492,-0.00829685808245906,-0.00454367128187516
"1807",-0.000531180416059707,-0.00639965808699117,-0.00429552812608569,-0.00683214464554072,0.00141664046019918,0.00108604050744132,-0.0036743459996581,-0.00931915146159878,0.000309931065455959,-0.00836828159099012
"1808",-0.0049428865682164,-0.00498645700951406,-0.0103538086391934,-0.0112098644499865,0.00264011690128263,0.000987071271906892,0.00545794903063279,-0.00651246414302431,0.00565318649217117,0.000383577422433889
"1809",0.000267187363282906,-0.00292351817172676,-0.00959006777714189,0.00206103867050556,0.00696041468430852,0.00394223699063834,0.00220080067376371,-0.00534084233235943,0.0146310949127437,-0.00268401243046767
"1810",-0.0112130585421767,-0.02157048165579,-0.0167251778264309,-0.0179993921395001,0.013450038259931,0.00589026793431291,-0.00322065532087623,-0.0126921226258663,0.0034153917507358,-0.00461366569400934
"1811",-0.00280808191849058,0.000856030068780989,-0.0116385028428202,0.00549871172457905,0.000184212167650522,0.0000975000288705452,0.000293594506176387,0.00074166343284765,0.00673170677617474,0.00540753876743816
"1812",0.00904355800433398,0.0130453541950233,0.01086969689379,0.0122396249363321,-0.00746366987304259,-0.00400121343534887,0.00161517715841319,0.0091403577866338,-0.0109692481907178,-0.0111410364454776
"1813",0.00713799248455071,0.00865526450420884,-0.000896090643081271,0.0138922608468424,0.00362076031693004,0.0024495165112095,0.00439722968435396,0.00538546160124698,-0.00774843518496227,0.00505051615747321
"1814",-0.00532891421618698,-0.0146504454250187,-0.00538126753103341,-0.0213140827423643,-0.00777058339206382,-0.00928545760997157,-0.0176590358026468,-0.0112005864164484,-0.019369155541615,-0.000386463282109228
"1815",0.00583963789758513,0.00127439146476638,-0.0144272567611762,0.00440748655482404,-0.00177146891699331,0.000197638831328728,0.00133713335543351,-0.0123123020782109,-0.00179557348100801,-0.00464046671164819
"1816",-0.00387839798110545,-0.00318194896424873,-0.00457483579759332,0.00619520481059088,0.0108341411660686,0.0018740911154953,0.00816026513760271,0.00170643626864408,0.0047708430723381,0.000777070152832904
"1817",-0.00413560471668872,0.000212873110862155,0.00367663335574586,0.00974860343881101,0.00711465639956321,0.000393850093857617,-0.0058863884568916,0.00325680982439525,-0.0178251808373535,-0.000388273345873769
"1818",0.00474579266067243,0.0129786616317988,0.00457882452032443,0.0114329634531083,-0.00376176751113144,-0.000590248662239334,0.00732220878428214,0.00998746970762032,0.0018228245363765,0.00660197167429399
"1819",-0.00719228514789438,-0.0018903071352383,0.00729271209442195,0.00226084906970514,0.00782763044631474,0.00423404150371143,-0.0111491180682278,-0.00494438716784373,-0.00791076630295806,-0.000771634106060737
"1820",-0.00210822719857107,0.00273568176848604,0.0144794790417586,0.0130324085868923,0.00502577796019121,0.000980561721375839,0.00481049497796104,0.00993760466733873,-0.0065386171265891,0.00888022757835838
"1821",0.00492998830236324,0.0062959344686595,0.0107046855690616,0.00791693673443739,-0.00563680770803188,-0.00352599234984241,0.00658283666982307,0.00984005650294084,-0.000240773745590395,0.000382775466384988
"1822",0.00819469244395821,0.00688197900710774,0,0.00662724017948402,-0.0024686954152493,0.0000977107317214898,0.00579679422268109,0.00292375962390978,-0.00762682253736069,-0.000765021771425012
"1823",0.00663031728726415,0.00683533661945801,0.00264783935353763,0.0117044323635678,-0.00854647812204168,-0.00206836289290824,0.00635461888311917,0.00218580275820734,-0.00177980744454487,-0.0122512563764504
"1824",0.00334678908861052,0.000411262927559219,0.00880299999772749,0.00192832216321759,-0.00574641835042611,-0.00434202845713816,0.000146618280187916,0.00799776128208207,0.00753708572442724,-0.00232554975998711
"1825",-0.00132374412424807,-0.00267323906349826,-0.00523572442126941,-0.00384911176026126,0.00438141198942166,0.00069356547034638,-0.00352355061232035,-0.00384701647810615,-0.00321751930501923,0.00815851687320612
"1826",-0.0118220608786495,-0.00371133677618907,-0.00438595952380005,-0.00265633413739375,0.00668303687203831,0.0061413609731229,0.00397803647325579,-0.000724194287114677,0.0133150583168988,0.00462429368806183
"1827",-0.0110514831843983,-0.00393207713491872,-0.0096916518707334,0.00435820754362815,0.0059925753349872,0.00236255167140587,0.00102732083779244,0.00458939106572487,-0.00525600063709475,-0.00230146453460378
"1828",0.00412313700769107,0.00332440386453148,-0.0213523263834662,0.0115720348688495,0.00238320514133727,0.00137477060966473,0.00557110099674474,0.0026447682026296,0.00944673734859536,0.0115339861699637
"1829",0.0107506979516336,0.0132532586991225,0.0145455469638154,0.00762637293761292,-0.00493735569678888,-0.000293815760705862,-0.000728892592357089,0.0115110996978012,0.00182412568242118,0.00266054900521828
"1830",-0.0210060175210964,-0.018393604400786,-0.0286737440150915,-0.0106434729064873,0.00928005538507892,0.00421846750274524,-0.00890004417704082,-0.0113801022067284,0.0054623337555415,0.000379147925316126
"1831",-0.00900828351083816,-0.00666265015781287,-0.00369009766495809,0,0.00810299977949569,0.00205137570704772,-0.00603562699812654,-0.00167822121833017,-0.000629887400521389,-0.00454719271475734
"1832",0.00787795809457204,0.00482099358022214,0.0138887688122635,-0.00215145287923191,-0.00261895822213198,-0.00155966085197978,0.00370262462309867,0.00384318706086728,0.00724807374143221,0.00913592825592224
"1833",0.00688768131216722,-0.00438055371047363,-0.000913175702619395,-0.0150933261259981,0.00624768986043733,0.00117177882899488,0.0106240341114714,0,-0.0184591320838347,0.000754344303005805
"1834",0.0104777701892877,0.0111040547812804,0.019195598090386,0.0126490188148054,0.00125939770902517,-0.00156010434966791,0.00598622342833655,0.00885396627770318,0.000398462035197555,0.0018846720080643
"1835",0.00139678399297871,0.00580191175218037,0.00269041209727328,0.00912777077247795,-0.0109639244821267,-0.00566605542585463,-0.00275748273610876,0.00450607327445107,-0.00629282295449407,0.00225738301863121
"1836",0.00348737036331603,0.00185408994464376,0,-0.00618881376029634,-0.000817753516185293,-0.000196425222284691,0.00422072864553913,-0.00283313704001498,-0.00408819238476954,-0.00337844807662935
"1837",0.00454454122985504,0.0065804469083568,-0.0071556322063655,-0.00263470125504828,0.00336483254536857,-0.000393192878138104,0.00333305165900533,0.00497267697827986,-0.00370250327917743,-0.000376565178978328
"1838",-0.00234201106975618,-0.00326881138606694,0.00270280367172582,-0.00720491760512521,0.00570983142981385,0.00255560912695874,-0.00303311391628747,-0.00282738654298265,-0.000161552756192895,-0.000753569186683123
"1839",0.00202732607207179,0.00143484398068439,-0.0035939255906694,0.000967756434502975,0.00189294983299537,-0.000294324814761326,0.00333235744291893,0.00307198388854935,0.00646409168610051,0.00603313866066468
"1840",-0.00819887516426732,-0.00450260180942419,-0.0063117824454112,-0.0135332251246404,0.00143938961055867,0.00137340169559952,-0.00346568969725458,-0.00494716314912969,0.00698460191047867,-0.00412292080413723
"1841",0.00316724708004945,0.0032892520362382,0.00544437450685731,0.00489972215719536,-0.00485067170326658,-0.0014687604725363,0.00521653224353757,0.00378807659942493,-0.00438493980706378,-0.00338731004097692
"1842",0.00465505656729226,0.00840173543987377,0.00270780628703293,0.00950744717367891,-0.00135379464749408,0.000882548128738447,0.000576546773165099,0.00589614314016562,-0.000160121720694795,0.00264346846756669
"1843",0.00298319666697355,0.00792519476467546,-0.00270049387274618,-0.00193174381837424,0.00415762850370394,0.00264582785171186,0.00446635130530693,0.0014067000607656,-0.00512574078867745,-0.00527299793137248
"1844",0.000105994845904123,0.00201623411358387,0.0126354296611935,0.00120968358850515,0.0107277264061754,0.00287913878123724,0.0077452485073668,0,-0.00338108192415798,-0.00757290238187724
"1845",-0.00143387481416746,-0.00321938729147464,-0.00178252425720637,0.00555822474261514,0.00615989311845055,0.00146462917687651,-0.000426865938578658,-0.000233681983857315,0.010177665343029,0.00267073913185523
"1846",0.00191442856884971,-0.000201915783506923,-0.00267837708684493,-0.00552750164620031,-0.00603348906177548,-0.000584837243926217,0.00355948240530513,-0.00117131576691465,0.0092755718739097,-0.00228319130765142
"1847",-0.0087038831478502,-0.00222075107647723,-0.0026858896702826,0.00459170791732766,0.00401745049850177,0.00117078611165433,-0.00368879057660321,0.00422061449153732,-0.00190142606638066,0.000762844652970829
"1848",0.00588912613728243,0.0036421497653143,-0.00448839880881946,0.00529243927383494,-0.00355644117168941,0.000779312293330836,0.0116776059915826,0.008171604036876,-0.0143673992451008,0.00266768573702603
"1849",-0.00106423382789622,0.000806686148989044,-0.00360664084886386,-0.00239314617251885,-0.00428275252276922,0.00107084568857951,0.00056313399288066,0.00115816855699036,0,-0.00304070567216974
"1850",0.00149151467943143,-0.00423063072143282,0.00814465104242279,-0.00167916334428819,-0.00322586705015238,-0.000777533947975195,-0.000140735021738725,0.00277571669359578,-0.000563743264294869,-0.00495612882897922
"1851",0.00973628152485961,0.00809228660531036,0.000897699483296099,0.0168190525559198,-0.00404509442043899,-0.0026286464643771,0.00211065446214875,0.00553609845933378,0.00676876723237352,0.00229889807629657
"1852",0.000895987788482433,-0.00220764431274112,0.0134527993805111,0.00378059999364488,0.00866459987145407,0.00390404992092863,-0.00589740971045716,0.00206473679032682,-0.00272133819879405,0.00458713250180853
"1853",-0.00473814246081894,-0.00140790958037917,-0.00530966526086762,0.00706223285339203,0.010828242421532,0.00456934410661902,0.00254252578854519,0.00251850342982185,0.00971107559728845,0.00456614763446561
"1854",-0.00878017875429915,-0.00382667472187925,-0.00978649921415009,-0.00935039246432579,0.00796678480165247,0.00358105880698179,-0.0016908123703776,-0.00159878015957249,-0.00826644159075485,-0.0060605625859117
"1855",0.00346858067329858,0.00141521399323219,0.0017970121434645,0.0132138960811725,-0.00280986893673851,-0.00212170902154707,0.00733863407993174,0.00365974959046911,-0.00216395773416589,0.00114331630053921
"1856",0.00366923952698639,-0.00141321399301375,0.00179381331322204,0,-0.00739827520947733,-0.00125687233397276,-0.00364227914235948,-0.000227919818463929,0.000642586345381391,-0.000761353473580639
"1857",-0.00630501477875878,-0.00545899969633479,-0.0116385028428202,-0.00815101214936065,0.00221810525326327,0.00290319305395759,-0.00309370826942146,-0.00934559287115533,0.000882966754166548,0.00190477512353748
"1858",0.0084244260113413,0.00833502510654527,0.0117755526457637,0.00774842799040232,-0.00610885419413365,-0.00154353721814848,-0.00394907008835532,0.00437172639439343,-0.0024059908187346,0.00190111471928089
"1859",0.00243210196587884,-0.00100806893090311,0.00984763109133535,0.00698994006076648,-0.00142519537560271,-0.00106325693732168,-0.000849645027694246,0.000916545835175198,0.0022509767847172,0.000759081054928057
"1860",0.00400842105743604,-0.000403653733504261,0.00975179569051798,-0.00185113527248593,0.00535242595027907,0.00203142237335285,0.0075112700656248,0.00595093153419479,-0.0012833560805865,0.00227528168495428
"1861",0.00614664609004456,0.00868145739238257,0.00790169725768242,-0.00857672582347957,0.00585591351496673,0.000289890446467433,0.00604864634911095,0.00227528698511881,-0.0213637776666328,-0.00832387743504726
"1862",-0.000730716839885348,-0.00460351756999255,-0.00435539536238472,0.00584528504516912,0.0123502976861689,0.00550079676455151,-0.00405489720966234,-0.0056752889549383,-0.0053344358692563,0.000381450015833007
"1863",0.00517273354774184,0.00361956622565396,0.0113734970373944,0.00278933292195349,-0.00531563259054024,-0.00124748862586277,0.00126354473830603,0.00525085306760498,-0.00214517332042496,0.000381422326485303
"1864",0.00161137141520729,0.00140262153968873,0.00173016833447481,-0.0136765568054023,-0.000438028700799342,-0.000769347923800123,0.00490738171853167,0.00272568927659123,-0.00421698355850864,-0.00762479245482162
"1865",0.00114193865585666,-0.00080036175319631,0.0120898332819503,0.00305531056989827,-0.00743376537852558,-0.00457565555563488,0.00181425046965655,0.00385050605333492,-0.00606163746574784,-0.00115257963929916
"1866",-0.000518269184423326,-0.0030036889722872,-0.00170636068428021,0.0056232684984252,-0.0123048305457399,-0.0050322912377474,-0.00125379179535812,-0.000677094836583514,0.00258984968896869,-0.000769141123897699
"1867",0.00202278296576086,-0.000803248259349187,0.00683732055956288,-0.00559182416972293,-0.000269377318871333,-0.000778307218645802,0.000976089738790709,-0.00293525049626331,-0.00208315970197215,-0.00269442259198116
"1868",0.00652189325267361,0.00824113086669098,0.00254680778650962,0.0105436150389238,0.000448232909567636,0.00146035908089082,0.0156034076184577,0.00407607873123239,0.00751504663468516,0.00115791773421514
"1869",0.00478284509750382,0.00737644661897896,0,0.00996989064181419,0,-0.000777777618001352,-0.00205761958654227,0.00902106831898686,-0.00041441238473694,0.00424041755856797
"1870",0.00102364660212606,-0.00178116556712116,-0.00084667857998999,0.00367308491620455,-0.00143361354409255,-0.00145868865856369,-0.0107218753328348,-0.00446997828625173,0.000331655747187964,0.00422274939862954
"1871",0.000102406309777203,-0.000792991725915848,-0.00847447252848188,0.0052607348007736,-0.00367960879265772,-0.0017537127871301,-0.00514072071779936,-0.00202042034285033,0.00613341887884933,-0.00267588302880972
"1872",-0.00347645803306362,-0.00674607502962132,0.00256400987983052,-0.00341299778662352,0.00180181907062948,0.00136609735753379,-0.00405043589402443,-0.00517446924216458,0.000164799408228111,-0.00268298369309872
"1873",-0.00707983246491317,0.000199723010386732,0.00341011622002529,-0.00479452939901115,0.00890098656586469,0.00389819280679315,-0.00294478230522977,-0.00271388399875871,0.0101309196892869,0.0142198340612605
"1874",0.00304833971058538,-0.00139799643712102,0.00509754528258166,0.000458901626537944,-0.000534651320851731,-0.00194148987271991,0.00253132305373938,-0.00385474796597296,0.00260926290451113,0
"1875",0.000824324895073225,0.000199891064859958,0,-0.00458636070616925,0.00249648418857085,0,-0.00505052930530037,-0.00455267686464456,-0.00439168025692638,0.00303140980953276
"1876",0.00277942521206631,0.000200018176093941,-0.00169058724820492,0.000230507637030586,-0.00791598030783702,-0.00418228391983666,0.00112835020585522,0.00114313166536162,-0.00114359583636003,0.00113334305133139
"1877",0.00733962940119692,0.00799674098325931,0.0135477641614032,0.011054864396834,0.00771056414396143,0.00527408345967428,0.00619715433978718,0.00776628592425488,0.00318939322202638,0.00415104216286699
"1878",0.00112084396847978,0.00238020317477372,0.0175439409543112,-0.0056945132873365,-0.0128118825310777,-0.00252601138897757,0.00769858841462145,0.00317333321235469,0.0348088698917237,0.00977074474588324
"1879",0.00203013690026754,-0.00257228293582024,0.000820890814442032,-0.00206206102419138,0.00757059949178363,0.00116850065981922,0.00347273923648328,0.00246976386921349,-0.00346622020692899,0.00186078579704874
"1880",-0.000305896005144413,-0.00178540564831142,-0.00820334653608379,-0.00206600690595715,-0.00313066420247776,-0.000680776221197887,-0.00235310976504843,-0.00547571804935576,0.00276678260869567,-0.0037147358734172
"1881",-0.00602429309365349,-0.00765393439722661,0,-0.000460273574217851,0.0101391796971788,0.00408912038965559,0.000461840606259756,-0.00183539243703978,0.00102487191209888,0.00149140393515124
"1882",0.00451971837642451,-0.00123382358825175,0.00349772104339041,0.00211110690924854,0.00257599730364122,0.00096990889415971,0,0.00666537971112735,0.0000787131813189124,0.00148918296182177
"1883",-0.000715804978160595,-0.00144146643328091,-0.00331949705915224,0.00115724464375511,0.00478382659237786,0.00261540985354336,-0.00111903321407636,0.00616431248825799,-0.00204736596657007,-0.00408908711055656
"1884",0.00194435735140219,0.00123732279764788,-0.00249796571444472,0.00231202379856321,-0.00149852479818791,0,0.00602068101256448,0.00476518735989995,-0.000552347497379868,-0.00186641921430597
"1885",-0.000510551348728905,0.00041196315535208,0.00500844234615272,-0.00276801834172646,0.00247253551976923,0.000773031873281926,-0.000834941038399539,-0.000903166594446003,0.0108952230887345,-0.00598361722093199
"1886",0.00669319919720501,0.00885311786498821,0.0174418048826614,0.00948407116817895,-0.00837249705347531,-0.0032691276607385,0.00250720961251516,0.00565082768785263,-0.00265538908612728,-0.00300977948909364
"1887",0.0010147407574066,0.00102041404391984,-0.00244887013351025,0.00595771776692477,-0.0106874541507177,-0.00407595422468021,-0.00111151898499928,0,0,-0.00188676673158761
"1888",0.00491841800236448,0.00550449090975391,-0.00327338408746769,0.00592271784440102,-0.00360097337953258,-0.00204643771171031,-0.00472952679881944,-0.0013483856798252,-0.0042286062074065,-0.00189041117318534
"1889",-0.00348156397277555,-0.0115571887087924,-0.00738923503891764,-0.000679144503998086,0.00731830828946256,0.00244138671429472,0.000978346633148552,-0.00472657545580646,-0.00110103016354102,-0.00795447621105305
"1890",-0.00642973826676296,-0.0133332208187137,-0.00330849196901972,-0.00453235231769167,0.0112118809452408,0.0045774224251629,0.00307174899760532,-0.00904575631799498,0.000393662424665209,-0.00267273931650935
"1891",0.00448407774949189,0.00395001069562029,0.00663897148264359,0.00569100265782074,0.000797995258442041,0.000193876771750423,0.00222721600672138,0.0088999662045377,0.00605962068151422,-0.00689125536772417
"1892",-0.00395704689147391,-0.0124249090370212,-0.0173124622299176,-0.00543251941109013,0.000266072598722467,0.00213248051463388,0.00319448126445931,0.000678707818244861,0.00547557119760866,0.00154199887714679
"1893",0.0013753525563851,-0.000629027368806767,0.00167788421560022,-0.00113775567874774,0.00637972009624965,0.00164488993895628,0.000692252283626349,-0.000452052745589016,0.00186716985428803,-0.00885304054897218
"1894",0.00503548742522919,0.00692404635446286,0.0117253555425232,0.00774682806027505,-0.00431434421083343,-0.00222121343364989,0.00456551591178234,0.00407034533344652,-0.02376143829602,0.00388352215418641
"1895",-0.00187288615920755,-0.00416755900240107,0.00331123053982019,-0.000678556874326164,-0.002033707183561,-0.000870909080377125,-0.000275383532566398,-0.000450393307190655,-0.00946549467494828,-0.00928428552675742
"1896",0.00370152342227126,0.0079513642783684,0.00165003871410008,0.00248881584433658,0.00531602966807543,0.00145248778018914,0.00371950390207676,0.00743581467549204,0.00353330124093221,0.00156178810632168
"1897",-0.0113659564376309,-0.0153621369460677,-0.00658975411046026,-0.0187318171084634,0.012603930186716,0.00580417564067415,-0.00590162045629383,-0.00849922868113939,0.0169640312317834,0.00233922971859379
"1898",0.0102192242763486,0.0078010540833946,0.00497521900899245,0.0156394965073616,-0.00322056674074533,-0.00201979288798404,0.00883593334866584,0.00924871094895896,-0.00755369447017684,-0.00661216291621969
"1899",-0.00187158354132888,-0.00460267278852278,-0.00165019624858609,0.00339677581567344,0.00497760199477604,0.000289184337599613,-0.00287388355626672,-0.00223518582848414,0.00166494097355763,0.00469848805988504
"1900",0.00435816040545078,0.00483385536418135,0.00330568999992309,0.00925290896180875,0.00208516752285459,0.0012524393446991,0.00425447866304385,0.00403205022430275,-0.00474907407785574,-0.00428688944394529
"1901",0.00221977984525501,0.00104610422793527,0.00082382879459475,0.000894465773663811,-0.00130091425287759,-0.0000958301681464047,0.00218712204443738,0.00401622067760199,-0.000954310497126021,0.00273980957205633
"1902",0.0000506538023961056,0.00522350119538406,-0.00493829782357291,0.0044681800235864,-0.0074663216038745,-0.00404199212584389,-0.00259113183145565,-0.00177764276329473,-0.010109894679751,-0.00117094414663099
"1903",-0.00468196256116626,-0.00706715897677701,0.00330851452979086,-0.00400349648938014,0.011808752978987,0.00386502079333417,-0.00560558822622703,-0.00823684561840987,0.011580241440776,0.00390772288067054
"1904",0.000404739677723143,-0.00167475924423599,0.00577092567972093,0.00692263799401638,-0.00138328812380106,-0.00115512811203589,0.00604934316557504,0.00157143365680579,-0.00166944111877387,-0.0019462560111887
"1905",-0.00429724662113629,-0.00293552603491976,-0.00245924165292732,-0.00598801913096558,0.00363651322210345,0.0013493175622914,-0.00464633484439936,-0.00112076523079463,-0.00302599931476344,-0.00312016237850077
"1906",0.00015246825083115,-0.0021029636909321,0.000821887677263433,-0.00490847213123313,-0.013887905840367,-0.00702475648994583,-0.000961219871999042,-0.000224064231017174,-0.00295523170020529,-0.00430358089483418
"1907",-0.0197482292051309,-0.0195996497209355,-0.0147784700778351,-0.0174886950420472,-0.00297409046526254,-0.000291145716284413,-0.0144313532731198,-0.0130162655907552,-0.0115357123842711,-0.0051080660694437
"1908",-0.0030555772445553,-0.0079536287255414,-0.000833076446691505,0.00547696893553695,0.00774082759736094,0.00588580367745517,-0.00195213788770787,-0.00250146576273846,0.0080233244835346,-0.00789890821798944
"1909",0.00722060548540204,0.00476693025359176,0.0016679060663003,0.00930569419662985,-0.00261845877299094,0.000579451708172973,0.00600820163525517,0.00364707841362133,-0.0031355443753549,0.00756371398691158
"1910",-0.0096961847274587,-0.011645133159359,-0.0158201315701111,-0.0152914239205459,0.00323801722467598,0.000482199922885007,-0.00888849833432814,-0.00885755170629499,-0.000967779675260627,-0.00474118489242559
"1911",0.000312606663197545,-0.00218226794395138,-0.0050762381848547,-0.00685084962680671,0.000610696609469441,0.000868131688249729,0.00182124304386333,-0.00779108535557671,0.0145313228094457,0.00635168079479187
"1912",-0.00541481575442437,-0.0113710968333004,-0.00340123968372119,-0.00390884412209436,0.00932879519211949,0.0045297434968441,0.00153877149627135,-0.00461869674690762,0.00405826377111906,0.00197235968110299
"1913",0.0115688735636004,0.00906896666684753,0.0017064237982003,0.00900261482141018,-0.00215973094372734,-0.000864045819085946,0.00754200454895604,0.00556871302251127,0.0000792677127912089,-0.00472426408615978
"1914",0.00289789737014901,0.00197260600031601,0.00936959838756724,0.0128119544500525,-0.0000865503237096332,-0.000479953383124676,0.00554478968595484,0.010844387775748,-0.00182267213213938,0.00158217528215698
"1915",-0.0013931989201853,-0.000437380893853034,-0.00168770376994021,0.00112909476556955,-0.00649304138414808,-0.00144121654726703,-0.00289500019922229,-0.000684997291881984,0.00023816291075085,-0.00631915096339819
"1916",0.00676920240443857,0.00415846271630604,0.00845324577846118,0.00541528309531736,0.0065354765035508,0.0032712604458125,0.0124430394427242,0.00799452492684583,0.00166679104161904,-0.000794901731337117
"1917",0.00472170202434929,0.00566698473985761,0.00167622598274431,0.00157090375237012,0.00805105217797752,0.00201354940425436,-0.000273373404978572,0.00702466804675672,0.000871640274286101,-0.011933134359741
"1918",-0.000204181176829077,-0.00130041769420364,0.00167367202697766,-0.00268873229909639,0.0109069327396443,0.00401901702544061,0.000956027830351758,0.00360017776443389,-0.00657109502923114,0.00402575128422056
"1919",0.00837941153136934,0.00781228760815122,0.00334175105868728,0.0096607390205754,-0.00993956118574923,-0.00314521717618821,0.0092798874616371,0.00470889566034627,-0.00414411848555662,-0.00842021728674447
"1920",0.00521852440255555,0.00193815117449025,0.0008327460823494,0.00467291229562505,-0.00308925187615983,-0.00105164953968584,0.000811187910631839,0.00490944822693185,-0.00224070904481988,0.00202189146360765
"1921",0.00267157523074668,-0.00429822713240768,-0.00582382774150259,-0.00199333676599356,-0.0016350155808269,-0.00296717934096213,0.00486331640620707,-0.00621767919305294,-0.00368943695861412,0.00282482003879458
"1922",0.00291587557172091,0.00561179104950815,0.00502101608093297,-0.00421684855678151,0.00560402555511663,0.00211187583706263,-0.000941006146704226,0.00335186174408619,-0.0107873449461653,0.00241449533829319
"1923",-0.00155391502775248,-0.0051514298842148,-0.00749380629913232,-0.00267414907226882,0.005572657369185,0.0000962106584510014,-0.00672860601097647,-0.00178229489545512,0.00252282721002994,-0.00160580016755862
"1924",0.00507025193930732,0.0101404129110128,0.00335585996131105,0.00737427459102014,0.00375158806545617,0.000766028402354513,-0.000406577767972482,0.00401622067760199,-0.00365292631458847,0.00160838290910359
"1925",0.000649374723376894,0.00170864165123286,-0.00501693094176303,0.00598934644011062,-0.00322757296307474,-0.000191443335700869,0,-0.0013332245486305,0.00496985505898406,0.000401439712543361
"1926",-0.000399298615902377,0.00405137459954186,-0.00420166901916208,0.00507174794738541,0.00852091072181516,0.00277634232509727,0.00162660314736862,0.00311535182444023,-0.000243194166894112,0.00160511449347278
"1927",-0.000549072221770253,-0.00594625195512721,-0.00253153263721062,-0.00987278233255318,0.00523876736653683,0.00133614797293835,-0.00094705108974491,-0.00510226444491235,0.00551410963347387,0.000801271114856617
"1928",0.00284774821510925,-0.000213725141077425,-0.00169198709048135,-0.00155108799133163,0.000672536410600166,0.0000953475271527893,0.00501139939866024,-0.00267560863317406,-0.00112902419354843,0.00200165638693472
"1929",-0.000498112630977432,-0.000854686019717943,0.0101693597294445,-0.00155367384194083,-0.0172503952320607,-0.00638817553887139,0.000538831336408307,-0.00268254450427619,-0.0178427174403138,-0.0143828316073027
"1930",-0.000548170686314964,0.00940976242690339,0.000839102285492999,0.0131142630852707,0.00556828265885656,0.00144146691969471,0.000269654390814056,0.0100873586050747,0.00411015200805331,0.00405353459188329
"1931",-0.00144623886341932,-0.00508475586135282,-0.00335304641240308,-0.00263279173491859,-0.0121825179228742,-0.00355093191972811,-0.00188535352247043,-0.00754534936834916,-0.00548505107678998,-0.00403716978450852
"1932",0.00449489647143952,0.00212958337661906,-0.00420529424557281,0.00857884833716338,-0.00189761759365159,0.000289108264018845,0.00944442354193242,0.00178901473182091,0.00477440719193911,-0.0016213804612808
"1933",-0.00258549436177857,-0.0131748600930298,-0.000844518537007954,-0.0117773519964512,0.000432272517926435,-0.00105942455676078,-0.00173753454122971,-0.0111606260257695,-0.0108962397328566,-0.00487208260272087
"1934",-0.00633109436096257,-0.000645683379021711,-0.00845308438217474,-0.0123593581622674,-0.000777318080501854,-0.00231299534584006,-0.00535561664407147,-0.0083522439802084,0.00115961232933959,-0.00815990734283745
"1935",0.00376254562324196,0.00409374800621021,0.0110827414644985,-0.00424585745595807,-0.00631026346458297,-0.00251183235306318,-0.0138644179946349,0.000455242722490201,-0.0050467525842619,-0.00699312305008326
"1936",0.00114959214249311,-0.00450638426465755,-0.00252955883876593,-0.00673239009688542,-0.00330543865203159,-0.00125949439616269,0.00122839972221667,-0.00750868779906855,-0.00656910848878922,-0.0049708498179174
"1937",-0.0058412126712688,-0.000646729906933152,-0.00338113691509812,-0.0106191708776778,-0.0104730255300668,-0.00378142143648863,-0.0287663753596186,-0.00320965745532442,-0.00912366276786081,-0.00791018072039307
"1938",-0.000753139455086482,0.000431423935869146,0.000848192432591155,-0.00502402893316722,0.00150001708534186,0.00184921391292692,-0.00407092945747656,-0.00850960870887763,0.00219633389583551,0.00125898658360835
"1939",0.00753811921723169,0.00366535919728372,0.00169485476286035,0.0130823872157899,-0.00405166835275983,-0.000291761977113558,0.00747048528915295,-0.0013915805247211,0.00160150877951359,0.00922045596687138
"1940",0.00134695098425497,-0.00386689228864101,-0.00846021236581751,-0.00928862354370485,-0.00256453120612554,-0.00252663346073234,-0.000699567622735486,-0.00627198697565379,-0.0108558527163871,-0.00415285260395082
"1941",0.00533010004812451,0.00927325161544856,0.00597271602382254,0.00137211221486,0.00319179218372434,-0.000682191114929176,-0.00727996869193215,0.0046753120124805,0.0020418410580072,-0.00959132395730922
"1942",-0.000901302307826368,-0.00491444461337853,0.00169629232584478,-0.00753604339975078,0.0127249150006634,0.00380256790600253,0.000563848904287623,-0.00503693483327516,-0.00585840555152328,-0.00294732818754173
"1943",-0.00772293098832855,-0.00365038000524232,-0.000846663704109685,-0.0151862199254711,0.00122229801984486,0.0021372648419149,-0.0088791123779226,-0.00329639499076406,-0.00204968834399821,-0.00844604763001489
"1944",-0.00572412045858006,-0.0129311841059101,-0.00169513214559902,-0.00560749437254637,0.00618786801494631,0.00213213408038881,-0.00568829813312155,-0.00685086612084151,0.00641848534734257,0
"1945",0.00782776184482348,0.00458520024430364,0.00594231895339914,0.0143325213403391,-0.00554376131420331,-0.00280493604835719,-0.00101042091137893,0.00404356031793962,-0.00467682831083038,0.00425901741067269
"1946",-0.0161355911841199,-0.0163007987438362,-0.00253153263721062,-0.0217743572428911,0.0118457201694837,0.00484964828649548,-0.00491179272958686,-0.0156363312737364,0.00290470731555637,-0.00212041208275215
"1947",0.00794543782139945,0.00419797135623634,0.00761419574445932,0.00449900713817653,-0.00146353709709679,-0.0021234465172878,0.0110336875100807,0.008905232846802,-0.00281115088858641,-0.0016999779678657
"1948",-0.00181900266699275,-0.00748077142131354,-0.00587752525454943,-0.0202730901268559,0.00801759590498441,0.00319255688221753,-0.000287150127015634,-0.0102575162776709,-0.000256270293119143,0.00595994531177846
"1949",-0.00263213212765268,-0.00066479761142757,-0.00591202139044567,0,-0.00564481587323529,-0.000868016315749065,-0.00603271355068846,-0.00192847509581673,-0.00700675046575028,-0.017350806458111
"1950",-0.0135523090612938,-0.0126444037218683,-0.0161428092882443,-0.0204524584507573,0.0193913522756126,0.00840152760914847,0.000577845379753583,-0.00748611481021955,0.00481884523551201,-0.0034453030602557
"1951",0.000154581627555883,-0.0112332875762298,-0.0189983744650919,0.0054041322478029,-0.0087120240044507,-0.00297225634507436,-0.00158844965317295,-0.00656917552345859,-0.000256906746345154,-0.00388940490539325
"1952",0.011009406426175,-0.00431709853715223,0.0123241789061004,0.00855111973629796,0.00426623099464063,-0.000288554209990521,0.00679859155642459,-0.000734789896899124,-0.0182456487621321,-0.00954442786635024
"1953",-0.00117046218171468,0.00821528186163212,-0.00260900574230316,0.01308149273586,0.000594837992746955,0.00163538774059901,0.00129304177781076,0.00171533094919663,0.0123898262595776,0.0127025911314935
"1954",-0.0154362826234513,-0.0212764866125663,-0.00610273246082693,-0.00884764106489955,0.0135008876574758,0.00585810861317659,-0.00588295398852023,-0.00831860512681448,0.00284410930659407,-0.00389276939652727
"1955",0.0174892487227372,0.0191950398663752,0.00614020448606012,0.0149577119382334,0.000251560517999794,0.00353234232861244,0.0190530267010709,0.0148038108537454,0.00953936052303739,-0.00390789288984161
"1956",-0.01983289685691,-0.0297254980282756,-0.0252832379605511,-0.0156878957724658,-0.00435561550192531,-0.0017123056757038,-0.00127493529722933,-0.0133721595471449,0.00144716096495134,-0.011769807888793
"1957",-0.011414468743304,-0.0137981096663137,-0.0143110060777361,-0.0217341413494089,0.00992671831662939,0.00390745065053588,-0.00141808779576336,-0.00566810510691929,-0.000425051006673338,-0.00352893522585584
"1958",-0.0164269664225847,-0.000236828188782345,-0.00907460538890459,0.0101209552165373,0.0060807467231947,0.00522094745310242,-0.00170421610793114,-0.00322162334630094,0.0079088445585116,0
"1959",0.00154750559342087,0.000711534914274559,0.00641020325195552,0.00586523369943781,0.00654076452852359,0.00198315326307164,0.0150803152581385,0.00273496925638406,0.00059060919483489,-0.0150509295657192
"1960",-0.00676641850973014,-0.0106659857711567,-0.00545933956403621,-0.0126337861023198,0.00789726948765246,0.00565525665574773,-0.00700773669548682,-0.00223166546435249,0.00337298265867214,-0.0125843292251807
"1961",-0.000858164131875117,-0.0103018829051812,-0.00365962155578181,-0.00910420412140578,-0.00636642363925077,-0.00271805327049068,0.00268185758675288,0.00447301304966663,0.00193296078549388,0.0100137531760711
"1962",0.01181085785087,0.0220284878889256,0.00459135451983972,0.0111744963115283,-0.0055851747305391,-0.00291331986491994,0.00506746299906924,0.00890678756056507,-0.00192923165635606,0.00360527101475738
"1963",0.00970974703059913,0.00450013079759226,0.0201097192056179,0.00294710418686539,0.00363463110398188,0.0014141523474438,0.0142856445232065,0.00882746442465576,0.00680733686540624,-0.00718459324177123
"1964",0.019810979382602,0.0150908475423022,-0.00179224618526275,0.00416259004664599,-0.00798327534701115,-0.00272948076722257,0.00952779714588381,0.0109383416441489,0.00183634386052556,0.00814114085177753
"1965",-0.0071109644482662,-0.011149955581254,0.000897683080043787,-0.00658364323271299,0.00107851571204742,-0.00028327337005829,-0.000410231412229733,-0.00769422367769668,-0.00566573085316779,-0.011215776547182
"1966",0.0116246955101691,0.0136248742155722,0.00627797453578949,-0.000245580449958371,-0.0088670049839461,-0.00415374920827349,0.00752611256532076,0.00993484998602057,-0.00687111636906701,0.0117966179513764
"1967",0.00769519922733619,0.00463491294362317,0.0035652273161817,0.00712021217747627,0.00100349519102227,0.000853110870947749,0.000407584241663317,0.0023993069271242,-0.00143434866944858,-0.00627794142929505
"1968",-0.00137448551612973,-0.00553634279152482,0.0017760627992589,-0.00780111539328465,0.00183766412326913,0.00104227767056098,0.00597299992823008,0.00191483191049158,-0.00245035914576019,-0.00270768346460881
"1969",0.0114701998672875,0.0153097563504263,0.00531924977536002,0.0201472143446881,-0.00625326266075621,-0.00246011417672698,0.00323899889067625,0.0102720894295376,0.000338810779922261,0.0081448253341041
"1970",-0.00151201309661309,-0.0105095361723544,0.00529084048421535,0.00144517353271412,0.00226539066753428,-0.0033197774058662,-0.00739860089922617,-0.00638426144402482,-0.0143098562965259,0.0116697308327325
"1971",0.00641060874582622,0.00600307398344357,0.0078948152321956,0.00937945823641995,0.000837059744207114,0.00104676035705875,0.00853780059306009,0.00975717070313076,-0.0104802161161337,-0.00842948025412049
"1972",0.0114352060364966,0.011935117708721,0.0496082740816859,0.00428892711083684,-0.00259296779418627,-0.00161617991975604,0.00752501805082795,0.0254533202529896,-0.0219636943838234,-0.00134235562090357
"1973",0.000545734924544572,-0.0131552322999143,0.00663346702706846,-0.00830372165874615,0.000000220853822563427,-0.000371812167010654,0.00773533450553643,-0.000919085797116526,-0.00452691267435068,-0.00896049769793583
"1974",-0.00346946931502468,-0.0022981222564501,-0.0263590164418407,0.000956759943795182,0.00310989000099315,-0.0000954039795244555,0.00119116310683665,-0.00897189819059874,0.000624155138222893,-0.0144666273901938
"1975",0.00631632067179555,0.00691086307739908,-0.0050762381848547,-0.0088428988374325,-0.00142421629287126,0.000286090859561217,0,-0.0078920481482343,-0.0216538939435582,0.0027524450020886
"1976",0.00400317744138623,-0.00388930849727853,-0.0127550894972008,-0.0122981667551652,-0.00646216758016482,-0.00305289638134887,-0.00422990299067161,-0.0138043633623181,0.000819710348668234,0.000914806340723828
"1977",0.000935337033453498,0.000229696544334912,-0.00344511282456128,0.00634763965603535,0.0114874835686027,0.00641164077427669,-0.000796658159103125,-0.0045076977784948,0.0281216243571611,0.00457041564431049
"1978",0.00314727453086672,0.00459252902501706,0.00777853083338353,0.00266871698111237,-0.00918565903995572,-0.00408874140939441,0.00451699513077086,0.00762637509452802,-0.0222183055482137,-0.00955414996961046
"1979",0.000980706043565593,0.00731415709877647,0.0060034745286035,-0.000967832146026248,0.000673996919088538,0.000095140524845716,-0.00251289225702067,0.00614944166303033,0.0143038386230658,0.0050528032285897
"1980",-0.00107750106515792,-0.0115724808682206,-0.00511502379857653,-0.00193775931158802,-0.000842294287337286,-0.000381416560663483,-0.00517103368794281,-0.00376121339467628,-0.00481971612977761,-0.00319922509623971
"1981",0.00112784297076796,0.00367295036406845,0.00856897870913009,-0.00266917226066077,0.0023606875571478,0.0016233042327003,0.00399862942844242,0.00283147287240926,0.00152464573991029,-0.0183402430648723
"1982",0.000244631829342756,-0.000914897227430878,0,0.00827251485384539,0.00487743542512731,0.00209768963127188,-0.00610648477720566,0.0070590121452796,0.0250739057056308,0.0107426411771041
"1983",0.000636409633649082,0.00228939078665213,-0.0161428092882443,-0.0106178684055914,-0.00251064805410406,-0.00114166470421917,0.00373975450159114,-0.00420584476571606,-0.00366906609881124,-0.00415900323180507
"1984",0.00577391128825355,0.0139333795269143,0.0138169525022147,0.00536601939606496,0.00276863812411254,0.00114296959226068,0.00479040176820678,0.00375428019184154,0.00876808394297024,-0.00510438663375412
"1985",-0.00160539522786218,0.000225402931300911,-0.00596247170117914,-0.000485056134431172,-0.00635884847055124,-0.00266405691786975,-0.00622466777291153,-0.00210376417342495,-0.0119078919102679,-0.00513052706809547
"1986",0.00175403868890167,-0.00427928264526023,-0.0102828071727715,-0.00169915367239226,0.00522034149429751,0.00181246782173194,0.00279859779867664,-0.00960413118094983,0.0103800228712174,0.00843884767950143
"1987",0.0053507362407843,0.00814281110142345,0.00779209560296468,0.0318502961058083,0.00603145610739508,0.00200019689950537,0.00730914710649899,0.00946065011700781,0.00461429562411375,0.0106925542322909
"1988",0.0028063591856784,0.00830153390517863,0.00171824579210078,-0.00824695380788465,0.00083253386196791,0.00114028844436698,0.00290246064600974,0.00163977279406002,-0.00242653611601129,-0.00873962635098224
"1989",-0.000723515050694123,0.00356055097155039,0.0025729477315386,-0.00641481865021021,0.00831936358721697,0.00246822039583439,0.00276229303978881,0.00233975834557487,0.00234554771657081,-0.00464030806755011
"1990",0.00255877233680879,0.00421265711627639,-0.00256634466086503,0.0126732029725345,0.00272308159737911,0.0017043884046728,0.00747737850413488,0.00210007600086715,-0.00190668231686641,-0.00233111440108369
"1991",-0.00211900669721377,-0.00684494091701304,-0.00343040983319887,-0.0200708331290741,0.00789936989492279,0.0038762599779536,0.00286454042934392,0.000465674216047374,-0.0264849157177869,-0.0457943004701402
"1992",-0.0069499276959557,-0.00111140509398056,0.00516342097096301,-0.0171083443732941,-0.00583412158846841,-0.00245284556788616,-0.00363548825305904,-0.000232587845821364,0.039871563287204,0.0205680919931677
"1993",0.00646403220779934,0.000222486954626788,0.00856154950503796,-0.000245168184261901,-0.00971212070544081,-0.00444411115873777,0.0035184617773063,0.00651929836889775,-0.0123520584602493,-0.0211132512505544
"1994",0.00386308743042552,-0.0017799134624652,-0.000848727395151183,0.0026974000931117,0.00390602136892393,0.000379663876195035,-0.000908938253656455,-0.000231446242199951,0.0103352701957204,-0.00588237341865872
"1995",-0.00110636090517113,-0.00401267154527041,-0.00254890121521767,0.00171192476020909,0.0083620049246409,0.0035127767748504,0.00155962479582583,-0.0115687671481495,-0.00386834859677898,-0.00295853949162506
"1996",0.00163722506435704,0.00492376536078987,0.000851897838427984,-0.00195326051061595,-0.0058292761769515,-0.00558209035300228,-0.00519081316722625,-0.0030428952870496,-0.012512918860362,-0.00247276535029672
"1997",-0.00668271879571203,-0.0075723037217138,-0.0161703782837974,-0.0146769862228523,0.0122223270520994,0.0033299360114365,0.00443534968590842,-0.0150271264957311,0.01179759678406,-0.0173525206683872
"1998",-0.000677571904304619,-0.00875217015864072,0.00519043372148431,-0.00943364527775714,0.00513999785317365,0.00369840952407796,0.0033766014354204,-0.00143018400341421,0.0208153655278578,0.0070634753146015
"1999",-0.0160315131282447,-0.0115463597796404,-0.0154904976458514,-0.0147873420213545,0.00730497443550338,0.00453560347369963,-0.00232957260520883,-0.00572937894600778,-0.00194604447168056,-0.0155310053935875
"2000",0.00507026624033147,-0.00366461783795857,0.00262206943970589,-0.00839478029956464,0.00411005985624291,-0.00169315740729181,0.000907937295734795,0.00432184385237244,-0.00228888608247602,-0.00916028487234122
"2001",-0.016161640013883,-0.0236781479490337,-0.00959015762875437,-0.0164187684095958,0.0135620462130273,0.00819675119546437,-0.0090734443822883,-0.0081281068454353,-0.00237911458273243,-0.00821792272696698
"2002",-0.00686955561528191,-0.0174241424673961,-0.019366062631066,-0.014345270716338,-0.00205878025213302,-0.00364442019180566,-0.0117723523047241,-0.0110872162903354,-0.0257218711959162,-0.0160538006646467
"2003",-0.00801962213510299,0.0119818576195743,0.000897683080043787,-0.00158769681022053,0.0123770170432866,0.00506441052257189,-0.00463267990034444,0.000974703919015329,0.00489551538504673,-0.00578939496770725
"2004",0.0196050283154798,0.0108925949826015,0.0167810092505662,0.0229868761841079,-0.00901252624908777,-0.00690548064517682,0.022340440885386,0.00998316446271152,-0.00591561563938092,0.00582310723543245
"2005",0.024728587356645,0.0210824267459637,0.0159715562718941,0.0136663449347862,-0.0177933044101736,-0.00563783018258313,0.0089750015350516,0.00867875640948168,0.00770110285379633,-0.00315774346202635
"2006",0.00425498596276563,-0.00145489773047092,0.00524015860263582,0.00700021654488769,0.0134458731534,0.00368571758632874,0.00206251584706152,0.0032046197392348,-0.00330008678592986,0.014783378020544
"2007",0.00460003159313627,0.00439409343622565,-0.00260650369137883,0.0139031947052812,0.0013504766948127,0,0.016467412831495,0.00816506444970178,-0.0193429821210155,-0.0182101106723288
"2008",0.00134947010554654,-0.00368411771420107,0.00174222595086215,-0.00914168820092831,-0.0198349464006992,-0.00828564773435092,-0.00506228229632322,-0.00119104058291286,0.0016880941353683,0.0100688091195851
"2009",0.0000962860091027196,0.00670225493450527,-0.00173919587866878,0.00230665789725082,0.00544276251695708,0.000722260145912257,-0.0041132807225307,0.00166927971934139,0.000266090123578033,-0.0131163498056155
"2010",0.00322475520766963,0.00114757910791696,0.00696869123317678,0.0079262412890484,0.00371145438728382,0.00133039538037494,0.00387207489806629,0.00428590199415524,0.0182673144879129,-0.00106324961847593
"2011",0.00134342992138947,-0.00802559290906424,-0.0103807556164052,-0.00608833118937402,0.007475019984168,0.00341547643148554,0.00437113137423695,-0.00379342886725387,-0.010101924408222,-0.00957959621759008
"2012",-0.00536611661158981,-0.00970863966936053,-0.0122376320452308,0.00204190388804948,0.00271308704361473,0.00113561149414543,-0.00102433368382504,-0.00309366920465648,0.0134600072747426,-0.00107467628639846
"2013",-0.00992303044702902,-0.00723642468045649,-0.00530981444047729,0.000764071730331661,0.00190943487565254,0.0011330370492082,-0.0153766965557564,-0.0076390627269971,-0.0140624569634321,-0.00753093793412274
"2014",-0.000535134801358805,-0.00493764159102039,0.00177954717979567,-0.013234718789659,0.0111178080018173,0.00509444748876908,0.0123634319445691,-0.00192437051203431,0.00440218340549059,-0.0119242345282613
"2015",-0.0180597103031903,-0.0300094745110773,-0.0115454375337561,-0.0177971678169465,0.0157087884401637,0.00610179379925335,0.00334273510285166,-0.00602553406286355,0.0150771473513824,-0.014262180473698
"2016",-0.00941873559958828,-0.0107186915624494,-0.0161724584748938,-0.00420200867257181,0.0180171201086141,0.00671790376131676,0.00730266204687502,-0.00339500017536021,0.01139896343526,-0.00946031160562877
"2017",0.0124609224601953,0.00935741754867925,0.0146118278230609,0.0216246857477227,-0.00197470104769104,-0.00018553819168543,0.01297375380923,0.0167885968555139,-0.00589141890646971,-0.00617957602536812
"2018",0.0177450797024776,0.0153694189426228,0.0126012224523444,0.0170365359545883,-0.0132429743758706,-0.00407836940594031,0.00565038727274025,0.0107681322824653,-0.00420852014085715,0.00395698354185292
"2019",-0.0080136126090472,-0.00624664408335973,-0.0106666351736541,-0.00329959107234123,0.0109526116754137,0.00493245419101407,0.000374443489223886,-0.000236786075058171,0.0113851990445886,-0.0016891660869599
"2020",-0.00783363719963259,0,-0.00359397710769649,-0.00814858394783557,0.0057217968314216,0.00351982450241617,0.00549216323532042,0.000947115857488967,0.0110864401997877,-0.0219966048061198
"2021",-0.00281269473890899,0.00435188256029839,0.0081155791555394,0.00872904070482861,0,0.00092311269976908,-0.00260719941121546,0.0082800534991645,-0.00337376861291772,-0.00403703159616031
"2022",-0.00603720162784405,-0.00192598066826988,-0.00178890329903403,-0.00559943657507245,0.00758636343875008,0.00461017355570381,0.00659636490168225,0.00375442320449193,-0.00160801450209835,0.0110017664138224
"2023",-0.00916038512425188,0.00603019941912497,0.0071683396517932,0.00230373477317025,0.0157354922720663,0.0085360068727951,0.00135992452856049,0.00186941037735622,0.0251759004392991,-0.0137458120305932
"2024",0.0131141482875423,0.0141449878274191,0.00889677096943875,0.00842685093101969,-0.0127493974509297,-0.00737175958305925,0.00851963355517871,0.017732284852978,0.0130642878606864,0.0191638030508074
"2025",0.00213264496779275,0.00732883347790247,0.00793675975594921,-0.00151952644154152,0.0132892881461804,0.00229198448184231,-0.00783512848443846,-0.00802355033246693,0.0137120473484831,-0.0136752043521947
"2026",0.00504817574570038,0.0077444153026458,0.00174968084698812,0.0220647638981257,-0.0115589848669275,-0.00475646293215759,-0.001481010331013,0.00762639584416647,0.000241594208734153,0.00635480048784021
"2027",0.0148706333356672,0.00302752425783304,0.00436678699512938,0.0191065386203737,-0.00359774126059598,-0.00248174677541391,0.0195256209263406,0.00366963700459122,0.00804958525196198,-0.00114808995632198
"2028",-0.00548273546784417,-0.00510782963597789,-0.00347832102381385,-0.00754805693555527,0.0139178868930414,0.00654218161839815,-0.00206080496185002,-0.000228195499267558,-0.00798530684376009,-0.00632181185090264
"2029",0.00234190865601502,0.0151690626418217,0.0113437588895577,0.000490461746892379,-0.00304204374139261,-0.0022886503859636,0.0098384334259205,0.00617140722626242,-0.00998152596035917,-0.0034702855386991
"2030",-0.0131906852038437,0.00137957328158023,0.001725807630784,-0.00539462843048311,0.00156314846740457,0.00137659415101377,-0.00132285536595234,-0.00477077145466476,0.0114643794042504,0.00522343606937192
"2031",-0.012824397559708,-0.0197429137632769,-0.001722834350116,-0.010847969600968,0.0163479960612152,0.0076960229442522,-0.00710581786432174,-0.0089021973498381,-0.00787784553251047,-0.0144341619889924
"2032",0.00924369399284086,0.0170959257994168,0.00862828952178196,0,-0.00658025223669656,-0.00354573538387559,0.00169819607328048,0.00967318101107573,-0.0215523905615361,-0.00468652079010523
"2033",-0.0125748422209055,-0.016117921963669,-0.0171087724435246,-0.0274178901285677,0.0177373004139467,0.00875992888184984,-0.0163480042706118,-0.0177920571524522,0.0222755461696662,0.0241318147701892
"2034",0.0123840047920647,0.0109993086848186,0.0104440220861803,0.0179395260554345,-0.00377554637404087,-0.00125033875630509,-0.0032008299642512,0.0188108386821693,-0.00834345099255041,0.0137930332837239
"2035",0.0144611710079967,0.0217591199891845,-0.001722834350116,0.0188821230173251,-0.0211661015412172,-0.00843722389575174,0.00926293555931279,0.00866200430184971,-0.0111909412055373,0.027777866916868
"2036",-0.00380768270708121,-0.0124601963479881,0.00517686141824858,-0.00494186361422544,0.00170891408957208,0.00164741040500016,-0.00293706142315775,-0.00949116709826847,0.00437834768166012,-0.0220628612013305
"2037",0.0100950098867001,0.0137644925479874,0.00858375901191244,0.00595971052168087,-0.0109794900670964,-0.00365389474762268,0.0104320027868503,0.0182519270423391,0.00172724951920977,0.0135363096736323
"2038",-0.00276542369034283,-0.015388165107001,-0.00851070516971408,-0.0170327408617651,-0.0177016174616804,-0.0111845657224664,-0.0263571328339789,-0.0100827927231709,-0.0258642086717776,0.00278243448269144
"2039",-0.00447564343949147,-0.00390690668763249,-0.0094418579493305,-0.00150682120969514,-0.00160354642716765,-0.0004638685305276,-0.00474071788910224,-0.014033552436324,0.00446728763037174,0.00998887909743806
"2040",0.0106530668110121,0.00945996239295699,0.0129982380264393,-0.0025151398247677,-0.00795408873833803,-0.00250370469904104,0.00350929932489796,0.00367300690801975,-0.00587393649196843,-0.0126373600584188
"2041",0.000580250730640275,-0.0061714303929048,0.0017107659101554,-0.00731211646461627,0.00185011398257262,-0.000372332538006392,-0.00212268774563895,-0.00251571271354911,-0.011817346063836,-0.00779065618397379
"2042",0.00961678992278148,0.0200091760730707,0.00683183985438274,0.0213361371581913,-0.00330870581042442,0.000372471221161463,0.010764579882248,0.00985989212039917,0.00230627829503716,0.015142982519029
"2043",0.00411654365028657,0.00338216798446345,0.0118744104346229,0.0114397018457635,-0.0102686287966286,-0.00334803268274897,-0.00544895129795797,0.00681212580995916,0.00545429539643072,0.0110495723323076
"2044",0.00157318926572714,0.00247198781758584,-0.000838299991074765,-0.00221277357763516,-0.015055884447902,-0.00709080195718259,-0.00286383725869743,-0.00270625741228858,-0.0166977534319948,0.000546553163430996
"2045",0.0000950460002353548,0.00403493628874996,0.0176174775830362,-0.00024622218170256,0.00594000723489341,0.0047923656677944,0.00849140259730863,0.0024872967035805,0.00284453059487055,-0.0120152404922721
"2046",-0.000713672634270801,-0.00178602376478154,0.00741976644898523,-0.00419050194060056,-0.00661385437011253,-0.00252477363123582,-0.0190687663729396,-0.00383483046540989,-0.00343814692928124,-0.00331676100198663
"2047",0.00600042773126064,0.0134197906654152,0.00900153103821011,0.00668301693785045,0.00293261777301357,-0.000562863228474098,0.00921513897787674,0.00543487949351085,-0.00569262539774673,-0.00388247916964912
"2048",-0.000142003414587366,-0.00441404520628019,-0.0056771160479181,-0.0100809660031115,0.0114588628834358,0.00459678202964642,0.00787931298873534,-0.00180174359375052,0.00130118842211302,-0.00668153796059567
"2049",0.00284063982317595,0.00620696940876031,0.00489388260914092,0.0144062850738247,0.0131262235553313,0.00662955610903238,-0.018862999361944,0.0051893439169417,-0.00147273672355541,0.000560530484758237
"2050",-0.000849622912622139,0.000660822878358447,-0.00243515663134941,-0.0019587982805821,0.00431842468959487,0.000928171623713503,0.0021502428475122,0.00246935211104771,0.00381741273959024,0.0151261328873129
"2051",-0.00118120717815828,-0.00462336620303561,0.00895050545415521,0.000245436661591603,-0.0136681722580416,-0.00593162652888191,-0.00845673101453304,-0.00335873216435389,0.00319795168188297,-0.00827820277748603
"2052",-0.00340637550809497,0.00176953376521083,-0.00403223478722536,-0.000735964721534255,0.00840810563746097,0.00354286441889284,0.00712875617220021,-0.00292060117853454,0.000775428620660046,0.0111296806566363
"2053",0.00631367672008953,0.00154556243316195,0.00242897764134797,-0.0014726841063768,-0.0186264287469354,-0.00744430413975694,0.00391795971725584,0.00856200976539689,-0.00413226569792469,-0.0143092756386252
"2054",-0.00410422528550325,-0.00859798237081355,-0.0048464249307113,-0.00762063971574189,-0.00362570267984419,-0.00215586857032457,-0.0026437096137526,-0.00513812448842488,-0.0018153440525589,0.00614179367706202
"2055",-0.00421564656494167,-0.00378014167592411,-0.00487004916024991,-0.0108990263800171,0.00031641523981385,0.00075147346248583,-0.00833165855859941,-0.00763533140855477,-0.00311769288024866,-0.00887895921922588
"2056",0.0010940025429873,0.00334829814943749,0.00570952971066463,-0.00150255818050582,-0.00126546665667493,0.000563500461968847,0.00330997243398712,-0.000452765123721388,-0.000955616358651601,-0.00391931914536592
"2057",-0.0140642092827504,-0.0180202306749787,-0.0016219671844836,-0.015299809276235,-0.0220917916347236,-0.0102270283367356,-0.0304491283936941,-0.0185645589943029,-0.0273043391304348,-0.0123666170244006
"2058",0.00414438220613156,0.00385143185130654,-0.00324929257765338,-0.00382055805893977,0.00923048844021723,0.00464500051491612,0.0088979088737553,-0.0129182755876219,0.000983372063442012,-0.00284572097699964
"2059",-0.0162216024812398,-0.0243735561314601,-0.01467005659221,-0.0222450628064117,0.0131578197560529,0.00424591199309332,-0.00492839989454252,-0.0170599681404072,-0.0049120567570593,-0.0131278504276504
"2060",-0.00234187494798022,0.000693840974329785,0.00909832210480599,0.00758376028738184,0.00728555587353164,0.00178527365328685,0.00143386967254711,0.00285318122457712,-0.00601326523089696,0.00520530925471774
"2061",0.0127137747982793,0.00809052416241274,0.022131248810545,0.00622896433584397,-0.000707305721271645,0.000937758549536039,0.0165297762349026,0.0109053764742246,-0.000270871331828459,-0.00460298819676297
"2062",-0.00613212194485546,-0.00710847078296961,0.00080191129730367,-0.0121228611083009,-0.00306851549848353,-0.00149884872104333,-0.00371307796835207,-0.00257940026424841,0.00144505056498345,-0.0202311155214705
"2063",0.0133603717539983,0.0145495878556592,0.00400649583883417,0.0120103981646256,0.00962749148428377,0.0034716252505167,0.0109240238890429,0.00940504026856992,-0.000631304129634969,-0.00118004618052503
"2064",-0.00297244076417358,-0.00409728934905795,0.00239423548439155,0.0116097593433102,0.00828516119189859,0.00205763754753452,-0.00089001738080341,-0.00652236081035007,-0.00541466483917807,-0.00708803408364778
"2065",0.0120214735467208,0.0237714287463384,0.0159236037298176,0.0244836451771657,0.0193027740128009,0.0114792354414828,0.0197224550331936,0.0192264615727302,0.0195989839361128,0.0273645963994336
"2066",-0.00456123602638814,-0.0136190820146114,-0.0117556082952225,-0.0169280595957948,-0.00509569680240463,-0.00470541445806394,-0.00149708234207591,-0.00253067111573513,-0.000711951569494884,-0.0167920756911898
"2067",0.00882682536420432,0.025124482865269,0.0158605308325934,0.0149405467650023,0.0052743455741564,0.00407840927101599,0.0242436644097497,0.019723197382328,0.0113990470086467,0.0135453445761553
"2068",-0.00194842340421686,0.00507837852622051,0.00468365679263694,0.00299406502695465,-0.00121670754258241,0.00129292158952055,-0.0014638233317833,0.00136207828715151,0.00633971119133592,0.0116211714476675
"2069",-0.00561916975341614,-0.00175758432813622,-0.00233098494621631,0.00398021618310218,0.00966877022035084,0.00304281524625871,-0.00806481294754069,0.00702796261621863,0.00244989935733742,-0.00804142308010869
"2070",-0.0146537445895898,-0.00528150308551967,-0.00233628331142288,-0.0158574703657881,-0.00844519049578352,-0.00432091958805891,-0.0165173558945306,-0.00562821233304256,0.00139655232608882,0.00289521423429195
"2071",-0.00238139059085585,-0.00973466473343387,-0.0101486180233251,-0.00931524263361239,-0.0155892498816956,-0.00563181817144365,-0.00568250096153633,-0.00950864525851158,0.00653708690306587,0.0121247840176284
"2072",0.00228940751492512,0.00178732411210825,0.00394338829669594,0.00279552035761177,0.0124372401575799,0.00389987225139432,0.00342887558894711,0.00571416157339977,-0.00363703662182968,-0.0199657933908359
"2073",0.0121998882476193,0.00356845078907764,0.00392779256698828,0.019259944430815,-0.00495955921006619,-0.0000926698250075519,0.0112644112136715,-0.00454547116177928,-0.011385346973498,0.0052385780379427
"2074",-0.00873929649605643,-0.0162223137567461,-0.0195617449638658,-0.00223775325402276,0.0021472916090195,0.00258985074702434,-0.00725901635031778,-0.010958944353794,-0.000791173626373598,-0.011580737745951
"2075",-0.00353627135417367,0.00880949559012811,0.00399031312850417,0.0124597238136683,0.0131343555001988,0.00475928032580408,-0.000126247430285886,0.00738688501490348,0.0170683963727469,0.0181605695309341
"2076",0.00359751507590667,0.00806094158694393,0.00874393633269754,0.0150134820614729,-0.0105954469730066,-0.00285102234062362,0.00668279547376294,0.00802024809712631,-0.00276815748733827,-0.00517835431905656
"2077",0.00673306568769316,0.00932906707252212,0.0118203712783425,0.0128517209441479,-0.00558374694750097,0.00129146504134536,0.0100199457584778,0.00727434653764125,0.0122311156508599,0.0127241223596799
"2078",-0.00264650739888017,-0.00154038441243065,0.0046729678501618,-0.0050277470170762,0.00838416778895579,0.000828992136571172,-0.0162449951393246,0.00157974712465947,-0.0049704429690558,0.00513984965216796
"2079",0.003377052287868,0.00110189934062377,0.00155029882825986,0.0209336990364595,0.000305594144071719,-0.000920374349456243,0.00277318915948155,0.00968910742730733,-0.00551201442156568,-0.0193180940344471
"2080",0.00442364057282485,0,0,0.00989850170284945,-0.0129646108918452,-0.00405359497685975,-0.0175990574195223,0.00290130444636683,-0.00692823238132634,0
"2081",0.00545696646833571,0.00330269491161306,0.00154798306794746,0.000700344466747715,0.00146803624108127,-0.000277586284879172,-0.000639700664318177,-0.000445261221740934,0.0113369061016291,0.0104287728250716
"2082",-0.00452267208123835,-0.0054860254841923,-0.00695508400084677,-0.00583049362825594,0.00138862368141268,0.00203541301188803,-0.00281674079142424,-0.0131344432663902,-0.0071570405522372,-0.00458721091733771
"2083",0.00191273984105633,0.00882616775625955,0.007003795990284,0.00445708496065711,0.00708805857217598,0.00295479041260061,0.002054197238744,0.00902329802950841,-0.00607952932151745,0.00460835039256935
"2084",0.00448706003062571,0.0050304387207758,0.00463700205435447,0.00700605231275575,-0.000841469476813628,0.000552870290872143,-0.0058942024724058,0.00268283238985689,0.00865080376353022,0.0200688264583102
"2085",-0.000284951710712744,0.00174103648727386,0.00230752860982797,0.00788496062188293,-0.00497687859430596,0.000735729114943462,0.0041243127465882,0.00312157170246063,-0.00346531231049119,0.0106800103349713
"2086",-0.011503677174857,-0.0134693184005579,-0.00767457416627282,-0.017487285969594,0.0114651927691065,0.00202276799016587,-0.00526268724973677,-0.0115582530505338,0.00495522042037044,-0.00222466379608099
"2087",0.00913690815330037,0.00110092859850752,0.00309365539145867,-0.000936802168555406,-0.00882470507040711,-0.00183517522507171,0.00129040684714909,-0.000674816315447191,-0.00761243092755071,-0.00445924791956631
"2088",-0.00119115681038551,0.00769916797536174,0.0154200692910731,0.00586014321106743,-0.00452826160259889,-0.00211412201295247,0.000773255625662994,-0.00224982982098676,0.0057531031576612,-0.00727885080943291
"2089",0.0049140585566938,0,0.00759307434636614,0.0107203858125371,-0.0152660119852167,-0.00580420038314367,0.00296215118884868,0.00270618935698641,-0.0134338277023877,0.00338416449252255
"2090",0.00251622263953699,0.00545728394425815,-0.000753587447927417,0.00737835576581269,0.00430625316579314,0.0030580395966151,0.00179740517453175,0.00202424646802557,0.00729159259788115,0.01236644346353
"2091",0.0023204914559174,0.00434219608023589,0.00377073795453886,0.00366206759027055,0.00623713791789982,0.00351052788893136,0.00166621545308132,0.00606071022415922,-0.0140415222731023,-0.000555353763433186
"2092",-0.00415787907645127,0.00713364159583807,-0.00225386632966174,0.00387684713195724,0,-0.00156529679387141,-0.00268694018577487,0.00178501275000653,0.0201680578460488,0
"2093",0.00317905315829314,0.000429218016660515,0.00301195723624259,0.00159013609525371,-0.0137911619444054,-0.00460980313622694,-0.000256594393970633,0.00289528111573811,0.0086707706811624,0.00166675834314023
"2094",-0.00411471937526375,-0.00836729975292516,-0.00900890062575699,-0.0124745004412555,-0.0122555788152973,-0.00370495616687894,-0.0196354836680002,-0.00644015135133535,-0.00704891245510331,0.00665542577805445
"2095",-0.0100205891438323,-0.00302897772813437,-0.0257577218186668,-0.0151582691432078,0.00174959712378264,-0.000279241290555343,-0.0116508787856126,-0.00916424698750617,-0.0176608169394716,0.00771362090786609
"2096",0.0108414445153988,0.00802949442495038,0.0124418748294668,0.00606337848240956,-0.0134611090124452,-0.00546681948143635,0.00529789970816763,0.00248124128214555,-0.00343702297138437,-0.0010934787598561
"2097",0.00284739391790878,-0.00172239476049219,0.00460819713843152,0.0057950171816985,-0.00943548209984535,-0.0020602946346816,0.00263527575814027,0.00607595238104497,0.0090201271839383,-0.000547337882276788
"2098",-0.011451721638971,-0.0148802219399641,-0.0191130812392187,-0.0108320408742525,-0.00138439954725744,-0.00168922649191539,-0.0219451007676443,-0.0136435649322304,0.00280455745494401,0.00821473346996493
"2099",-0.00411688146435385,0.00678644927041216,-0.000779410230338451,-0.0123484900106433,-0.0171204766595336,-0.00488831738712492,-0.00268688571266462,-0.00680282074485217,-0.000524357638950534,0
"2100",0.00398971060180497,-0.00413152139034834,0.00155988831780851,-0.00141546636965351,0.0134374424027568,0.00425114810045346,0.0132024050990676,-0.00639268719026087,-0.00821968338387813,-0.0157523714176044
"2101",0.0131660941726204,0.024890911388797,0.0233645013751749,0.012756832060153,0.00270103986904879,0.00385655478491209,0.0152901608730895,0.0238970853255613,0.00484925947538795,0.00551868825165203
"2102",-0.00477272836221998,-0.00447384949530361,-0.0159816979883729,-0.00956373500641206,-0.0243245865889097,-0.00983915153085058,-0.0145364481688911,-0.00897660385715893,-0.00386068260190675,-0.00439071958871129
"2103",-0.00299131612741299,-0.0038517847726014,0,-0.00329730129810679,0.00259329470989411,0.000757205439993802,0.0029234858768119,-0.00181169099839285,0.00854400606486383,0.01047394718828
"2104",0.000190480128019033,0.00644467064314336,0.00618714302101031,0.00189050733921015,-0.00801054693144443,-0.00132388583180931,-0.00834733962444023,0.0111162913568572,0.0179039563318777,0.00109120500779669
"2105",0.0104275612338232,0.0164353307568916,0.00538053340948474,0.00990561105712007,0.0026915991508365,0.00340908386580896,0.0181719996765111,0.00964768235812219,0.00540537952624498,0.00599463697079994
"2106",0.00108382677576735,-0.00146984266137973,0.00458707979572326,0.0077067829123596,0.0200506748705891,0.0071715422916645,0.0082678757059671,0.00866639511408596,0.00298684929168802,-0.000541704379498187
"2107",0.00310682970910703,-0.00546800683090543,0.00837151497176469,-0.0101971494510703,-0.0167778927380077,-0.00674590810341835,-0.00299364010303771,-0.00837152514099149,-0.0000851016768919077,-0.00271010147902528
"2108",-0.00032853496693741,-0.00338330770521023,0.00075462255427583,0.00163909210715674,-0.00886647493902049,-0.00443358033830854,-0.00130552571069231,-0.000888664985084553,-0.0138699629136307,-0.0211955866319149
"2109",-0.000704154091032083,0.00297037068408623,0,-0.000701281173385859,0.00168781731071599,0.00217922325395414,-0.00209156858695658,-0.000444609467145973,0.00163951161998011,-0.00222107217221601
"2110",0.00291228937319521,0.00571189427984109,0.00377073795453886,-0.00350876192432548,0.013986133559744,0.00595660928645447,-0.00458486334718,0.000222122672990821,-0.00335975183735771,0.0122427460883201
"2111",-0.00238849054143142,-0.0094656106981601,-0.00225386632966174,0.00328628106035844,0.000415430700419606,-0.00225586457115767,0.000262988665556518,-0.00556028963142174,-0.000777975611064519,-0.010995183959485
"2112",-0.0107518591470216,-0.0205988827420454,-0.0128012368139586,-0.0159100791406158,0.0171093513794323,0.00621729364177392,-0.00605155686584391,-0.0138671178278663,-0.014619325512445,-0.0194552740661222
"2113",0.00949222266537042,0.012575898331286,0.00686504000384036,0.000237584735121033,0.0022868036135657,-0.000561653428597819,0.0075448579383961,0.00249450594840939,-0.000175621098213563,-0.0136053739085655
"2114",-0.00112810465237523,0.00064228581169834,-0.00227287428307532,-0.0130733876055154,-0.00244440682415537,0.000936350612388503,-0.000657124450384128,-0.00610837268345477,0.00114143472773232,0.00517234311863457
"2115",-0.00621307828379081,-0.0113416352799512,-0.0091115903927883,-0.00963385817036455,0.00220541497723725,0.000561443352620428,-0.0107796085098693,-0.0102433719211309,0.000701640081607779,0.0125786219037087
"2116",0.00203664436815076,-0.00692643524608527,0.00459777055074828,-0.00389113768139526,-0.010747739074507,-0.00441201089310195,0.00970137912355584,0.00183977983909855,-0.000876406676185937,-0.00225858023963132
"2117",-0.00099282115181909,0.0076286112337911,-0.00228833287973562,0.00390633777952543,-0.0139519305637988,-0.0069628541706811,-0.00816031769877568,-0.00114782326774754,0.00403507894736843,0.0118846210882944
"2118",0.00264954073581558,0.0086523320742502,0.00382262868569572,-0.0051070060142564,-0.0160748825384622,-0.00852730327087325,-0.0120751177393947,-0.00459678298209887,-0.00716407484854154,-0.0128636462591393
"2119",-0.00844647853750868,-0.0113660564118058,-0.006854521053545,-0.0151552914977839,0.0130188812696757,0.00487333167951221,-0.000940794838816594,-0.00923592987427313,-0.00703980118831227,-0.00906514926579005
"2120",-0.00171332875106378,-0.0140997859321327,-0.00613509612626495,-0.00446750892255421,-0.0121799449890934,-0.00722752883780298,-0.0120994239377238,-0.0146814458924173,-0.0053172458460562,0.00457409782496465
"2121",-0.00614943198803963,-0.000439983915517028,-0.00540114552153914,-0.000249330415946214,-0.00110531255402013,0.00143687914970814,-0.00204144651770466,-0.00402108678724866,0.00294014616785709,0.000569144195399662
"2122",-0.000144372960119599,-0.00506272835546406,-0.0100852123687302,-0.00598486453006397,-0.00791682151674622,-0.00325240287721684,-0.00722770417122043,0.00522441580692923,0.00222084036599446,0.015927265450697
"2123",0.0119936399927618,0.025000134727625,0.0164576178674962,0.01455073923432,-0.00875238208509166,-0.0038387562162534,0.00714278654826805,0.0181906094216553,0.00850912072327614,0.0039193191453657
"2124",0.00322349770211305,0.00215810858299492,0.00462596225174328,-0.00494561234091917,0.0210352014333548,0.0079001427459473,0.0079104009831954,0.00255192781875824,-0.00457019691132188,-0.00892358463847098
"2125",-0.00765474281905421,-0.00969190554299504,-0.00537227474894364,0,0,-0.000573838627972778,-0.00189415887822275,-0.00485976604704164,-0.000264868439610377,-0.010129466925154
"2126",-0.00428565340434983,-0.010874289796337,0.0030866408515231,-0.0111829550693209,0.00161113728340312,0.00239092268763441,-0.00515200230267598,-0.000697792826756416,0.00441579075114928,-0.00454797665417239
"2127",0.00545172979287112,0.00065961669279524,-0.00461559950994483,0.000251419932364216,0.00787177851241938,0.0038164145776125,0.00844920954922634,0.000232481606111001,-0.00360505573889769,0.00285547202898218
"2128",0.00161707550326584,-0.00131836377083994,-0.00850059070470233,0.00603031365049445,-0.00772647812874372,0.000570537344617872,0.00621623760420564,-0.0030243729148981,0.00467700317684439,0.00284745874768899
"2129",0.0103994164054775,0.0127612099694838,0.000779262294557048,0.00924065356865778,-0.00490884408931846,-0.000760310514036022,0.0138329611954167,0.00560095377468128,0.0129117437489985,0
"2130",-0.0044393111880372,-0.00391048611150291,0.000778887807170614,-0.00866133601621433,0.012842925352923,0.00532401991577003,-0.00649098994341823,-0.00359023653346646,-0.00173427852930974,-0.00908585572589227
"2131",0.00512320815705247,0.0233370562562201,0.0155641552067913,0.0144782371381589,-0.0204061246450059,-0.00841615123695394,-0.00986654354203165,0.0101269592149413,-0.0128561845155615,0.00343846653051139
"2132",0.000707992962514892,-0.00149186957653658,0.0114943744333482,0.00984276822675856,-0.00600094430706521,-0.00305170901455509,-0.00484811692387255,0.00373050737714009,-0.00659978886483448,0.0119930413004823
"2133",-0.00726290161408316,-0.00787786230800114,-0.010606109874057,-0.0070664575880921,0.00862434152864666,0.0029654162638697,-0.00562481002717929,-0.00766542229949407,-0.00265748075699779,-0.00677197507159488
"2134",-0.00304033167630813,0,0.00200097246859188,-0.00343618807021773,-0.00350562246188768,-0.00247966095453778,-0.0094742630682263,0.000701976572409002,-0.00133221427594676,0.00113634815293406
"2135",-0.000190782644676757,0,0.00460821940299394,-0.00942719890863131,-0.0112408230035713,-0.00478063053157674,0.00485166048642283,0.000233766547662606,0.00106720026561358,0.00454040856141935
"2136",-0.0209700528299418,-0.0335599562343512,-0.0252293793219545,-0.0222889887433528,0.0264687674216355,0.0116247277700927,-0.0160022777326081,-0.0240876373560918,0.00453093469315813,-0.00451988643037415
"2137",0.00209318502478051,-0.00748970449930952,0.00470597495388425,0.0148566199005866,-0.00693275860754616,-0.00275420837496609,-0.000420581851782509,0.00311519875064414,-0.00619082869019183,0.0215664003574805
"2138",0.00801532764409907,0.00548814370178352,0.00702564601085265,-0.000757168457274915,-0.0134979403943855,-0.00522636965864054,0.0152874362684248,0.00334460659300873,-0.00347067713435945,-0.0122220558958132
"2139",-0.000915606377680733,-0.0002275189398252,0,0.00479907129402646,0.00328637241120822,0.00354726480066714,0.00221047234394089,-0.00214290789320903,-0.00196464541977193,-0.00168738161556348
"2140",-0.00284574464036014,-0.0245677463598537,-0.00697663067339305,-0.0279034200011654,0.0185347542728374,0.00706992387834093,0.00454833881004846,-0.00978264367666826,0.00268428771144791,-0.0326760730635546
"2141",0.0062886938481177,-0.000932681593462714,0.00234179776477283,-0.0149986837493136,0.00939502551941129,0.00265612637924129,0.0153678479848511,0.00192763297168796,-0.0116008925861304,-0.00582415211058229
"2142",-0.0167774689501847,-0.014706065428325,-0.0412771615979164,-0.0343921973992904,0.0086365218712805,0.00397371291625426,-0.00527027224867949,-0.0264551375289911,0.00297936072626648,-0.00468652079010523
"2143",0.00180915428887074,0.0175313362515475,0.0121852131180118,0.0193040493718217,-0.0197023265598012,-0.00697327815946658,-0.00475472397400589,0.00963434505717808,0.00243050688380619,0.0117715903659563
"2144",0.0125913978388434,0.0419091522691211,0.0160512172206979,0.0253398085420107,-0.0158581877632955,-0.00692829238612869,0.00696164458762993,0.020063413641733,0.00116735810733348,0.00465380499809842
"2145",0.0110372680855471,0.000670533341460944,0.0134282716684846,0.00676401917808733,-0.00310229048062682,-0.00267599667476548,0.00149098015538973,0.0115137544714301,-0.00448470722907357,0.000579150118952709
"2146",0.00433818192022994,0.00848599470016631,0.00623529077560958,0.00180870689289936,0.00328453918396709,0.00316214817917326,0.00270682688082813,0.00758840224891322,-0.00225245521673045,-0.00347241290050826
"2147",-0.000332292180052485,-0.00465019110832954,-0.00077459466577845,-0.0113489999819608,0.0105970061697793,0.00382080264825735,0.000945072964895655,-0.00282440516245208,-0.00523743914100483,-0.0116142449742631
"2148",0.00802427657181659,0.00912127424723441,0.00387591290059119,0.0125229096246389,0.00690555682634542,-0.000380417251551357,0.00714773083733156,0.00991295217954646,-0.00363110008601675,-0.00470034876032666
"2149",0.000847952883457737,-0.00352725277059718,0.00231666891479132,-0.00128833305720744,0.00516461015027181,0.0000953466920246004,-0.00388334445663918,0.000467372410373201,-0.0101129735766586,-0.0053127963211177
"2150",0.000517519192555271,0.00309728355771499,0,-0.00645000364314752,-0.00421154133988899,-0.00199925028505765,0.00174780982258138,-0.00186883125469273,-0.0271514491090392,-0.0160238240596492
"2151",-0.00395116915285032,-0.0037495277127978,-0.00308171091841491,0.000259731551730535,0.00541351235212084,0.00276574768053961,-0.00362337662733181,-0.00397850581154902,-0.00312198684357579,0.00422195857957752
"2152",-0.00179469737313753,-0.00730575441686443,-0.00463670988986586,-0.014278499929954,0.00622545533416319,0.00123662100492061,0.00282829265599482,-0.00258442484879207,-0.00540950919399696,-0.0144144029424824
"2153",-0.00562987191849795,-0.00289917244495264,-0.000776482597506956,-0.00974451885067695,0.0124585698953876,0.00408462061588577,-0.00711803657292698,-0.0110721967541599,-0.0044847422380323,-0.00853139209343812
"2154",-0.0103718175535955,-0.0118540602973378,-0.00932394189529828,-0.0143614983129285,0.00247750081138642,0.000946597432893048,0.000270575613710022,-0.00262031991282485,0.00977663165385545,-0.00799018329028789
"2155",-0.00581773366541882,-0.00792233822888477,-0.0039215964243291,-0.0188885465042907,0.00535453198061075,0.00330771362374582,0.00216364787610845,-0.00286572678798669,-0.00465113440248954,-0.0192069322486307
"2156",0.0122832732101361,0.0134612263637814,0.00472458751465887,0.010176214688481,-0.00729242030562671,-0.00282607958064551,0.00188912266667729,0.0124551716719983,0.0015258058218024,0.00821227311896955
"2157",0.00687891870183699,0.00225132475439871,0.00391843791884727,0.00980117236630584,-0.00371468824530008,-0.00141731903456188,0.00511795942349491,0,0.0014283089343452,0.00313291822478545
"2158",0.000237491753570129,-0.000224708155990405,0.00156126168898196,-0.00997571723645219,0.00770515323650156,0.0011355475479875,-0.00375198307375868,-0.00260252849842257,-0.00855758312365851,-0.00374779901424127
"2159",-0.00151805896858048,0.00629069855297137,0.0077941187262327,0.0108932015964092,0.00739956918181672,0.00585883130350706,0.00645608664849928,0.00308342637742687,0.00632974987042534,-0.013793109233514
"2160",-0.00337299162336402,0.000223252488680048,-0.00386692012852963,-0.0167024781986888,0.0105264767407549,0.00304862119241123,0.00494444587662102,-0.00425571214456955,-0.00791005432192893,-0.0165288315302095
"2161",-0.00195400070448593,-0.00267853299718046,-0.00155286046872471,0.0035616282617299,-0.00793193206334464,-0.00515966119892997,-0.00518612463555013,0.00403645650821849,0.00201729110503912,0.00581769849731795
"2162",0.00329518431833442,0.00671436769818978,0.00622082966701987,0.000272849882013482,-0.0075059767232335,-0.00386580941105386,-0.00427754955643334,0.00496708890073028,-0.00364296814577625,-0.00385605447913029
"2163",-0.00818765294286794,-0.00111162278171673,-0.00309115382533776,-0.00873348050422051,0.00887758746754796,0.00350239860248203,0,-0.00117691283141264,0.00442604637736932,-0.00064521886644664
"2164",-0.00192006441156345,-0.0040063257456594,0.00310073868558702,-0.000550693664033597,0.0131184908276887,0.00396208002590592,0.00349020502795816,-0.000942453818183364,0.00249068878715097,-0.0038734139922495
"2165",0.0125993416484562,0.0118437442743728,0.0146832621202542,0.0168044786335639,-0.012385128921667,-0.00413443642998934,0.000134099342269156,0.00778305929077083,0.0102245482995786,0.0213869496870762
"2166",-0.00902297383022821,-0.0136925657757676,-0.0175172062151208,-0.0219454836760518,0.0158790187005693,0.00660420358998692,0.00668788311428492,-0.0142757226756955,0.00510784141971388,-0.0133249515791739
"2167",0.00119780130100677,-0.00582186648346783,-0.00620145645838888,-0.0155123178519413,-0.00545058903448115,-0.000374535267901321,0.00146176364858452,-0.00261179717225668,0.0140221905887035,-0.00321539024234307
"2168",-0.00124447989707266,-0.00292787753730828,0.00780011421873894,-0.00168812077928804,-0.00322410333911094,-0.00262526521168605,0.00199018845648857,0.00166666108620017,-0.0082598515081207,-0.00451613365891079
"2169",0.00364238627869584,0.00158122616145739,0,0.00140893753250326,0.00234494719749856,-0.00103421264879622,0.00569370104280686,0.00617835669189049,-0.0000936084587908059,-0.00648092618506435
"2170",0.00558678301452931,-0.00360839399780821,0.00232202740308063,-0.0109765315932372,0.00451753364525076,0.00178768364830617,0.00750513677595332,-0.000235937097971206,0.00262048671259696,-0.00391384098282155
"2171",-0.00289655761971896,-0.005658886248044,-0.00694977759190962,-0.010814060135763,-0.00787028781362742,-0.00159676255920504,0.00078398644620048,-0.00519684108186136,-0.000186651736768018,-0.00523909389894606
"2172",-0.00790554701329149,-0.00956068315264735,-0.0108863208058256,-0.0123703406666167,0.00987564542687114,0.00611579529221329,-0.00548446391686519,-0.00474991273787839,0.0134441414112207,-0.0111914887418054
"2173",-0.0208811604169064,-0.0216042511988987,-0.0298743461908856,-0.0157296202873517,0.0100992218562976,0.00271199940023714,-0.00774667146103403,-0.0174184048842674,0.0174113214902445,0.00266307934858157
"2174",-0.0301028023021378,-0.021611324966379,-0.0340356933225653,-0.030778334802554,0.00301578417445625,0.00401054891812147,-0.0195847288344548,-0.0206410874571306,0.006247690940824,-0.0166002437314864
"2175",-0.0421067909287234,-0.0268907692789102,-0.0352348257364755,-0.0436640344914877,-0.00031686608868986,0.00167233124466715,-0.046699961667269,-0.0453754190156463,-0.00539906430484294,-0.0249831944517125
"2176",-0.0117674819728253,0.00616817270045433,0.00608687296800836,0.0127713028135317,-0.0160650477467194,-0.00547161355290193,-0.0252018269398729,0.0070127770687336,-0.0123947798099592,0.00415521063827451
"2177",0.0383936027431702,0.0166747790970849,0.0397580652682827,0.0331021777847089,-0.0193035166699025,-0.00615445544295645,0.0249817950808431,0.0201186983604777,-0.0136497429956122,-0.00620695348291322
"2178",0.0247352459916323,0.0108541181514457,0.0182876006150599,0.0442478364765475,0.000573934578958601,-0.000562968137750031,0.0201218699957466,0.0199746993634025,0.000557304737759834,0.0360860590358638
"2179",0.0000501048404741855,-0.00238615697177935,0.00489805568691937,-0.0128580632065616,0.00295108335615302,0.000187453353823752,-0.00111112014456327,-0.0101636049585033,0.00900393551460321,0.0261219592799926
"2180",-0.00807917318208962,-0.00454442849140002,-0.0154347187023525,0.00177604208841475,-0.00768223845022142,-0.001689282089954,-0.0198860542184029,-0.0120211472317938,0.00110398347113105,0.0241513737615482
"2181",-0.0298477649326073,-0.0285920857338701,-0.0453795722233137,-0.0387112607481843,0.00720536281378314,0.00449171904836665,-0.0190124517914777,-0.0263622627305049,0.00349197757765118,-0.0331421357263799
"2182",0.018981245494792,0.0140984930958568,0.018150584318078,0.0144479868310672,-0.00860430052906469,-0.00271864572880764,0.0107030629845959,0.0179637898568914,-0.00531130051221518,0.00856963182897941
"2183",0.000716354006460751,0.00146344896062267,0.00763994257779532,0.0039394779177504,0.00487655323052705,0.00244417293362131,0.00200315065783085,-0.00306901515148461,-0.00718106222110859,0.00653585802039114
"2184",-0.01513673849902,-0.0211883942115232,-0.0320135339286063,-0.0298823055565421,0.00913053278984099,0.00309453732483078,-0.018994318526194,-0.0218057514870087,-0.00324553053581345,-0.012337627793219
"2185",0.025131038236041,0.0291116653825398,0.0234987124174919,0.0317360797201094,-0.014753735426546,-0.0043937523424219,0.0151405726238329,0.0251767353680699,0.000279086431837161,0.00723212063576195
"2186",-0.0133716684641875,-0.00531920019536269,-0.00170056853691969,-0.00512651303208156,0.00479833078366609,0.000375476521343066,-0.0121900527807146,-0.013814268453044,-0.0129278277416619,-0.0130548529148178
"2187",0.00544152356088112,0.00947979923058706,-0.000851767166973549,0.0103061956902502,-0.00675157542637894,-0.0022522906184409,0.00116154830146931,0.00985762418203384,0.00235560168724014,0.00859783403115144
"2188",0.00454447370921107,-0.000963027235667768,0.000852493292770262,0.00390040588815266,0.00630015228408087,0.00263370173699373,0.0163860547558181,0.0020545837014756,-0.00206799216209796,-0.00131145753062911
"2189",-0.00371056427080063,-0.0106050666656551,-0.00255541639653756,-0.00149452669328987,0.0015655342129155,0.000938130395796044,-0.000570645776742373,-0.00281954662348094,0.000565156346452156,-0.0124754099800847
"2190",0.0124993451787259,0.00682103617884944,0.00768582072454271,0.00957801140366032,-0.0191646552486338,-0.00787382571002815,0.00842273908504287,0.00385600872698966,-0.00301260588389562,0.00332449124458023
"2191",0.00866654543069179,0.0164529582078587,0.00847436121075895,0.0243107063171968,-0.00377338177146158,-0.000283239495014298,0.012882145342666,0.00717032648609428,0.0133144095691329,0.0165673099142225
"2192",-0.00224798474247956,0.00285652931903368,-0.000840246977840353,-0.00231530176439187,0.0122052632270604,0.00831647803017099,0.00978360273777001,0.00101711147160688,0.0102507317165359,-0.00651901687994838
"2193",-0.0163412234823096,-0.0256351051861363,-0.0319596169840316,-0.0185670411035254,0.0153844411139754,0.00468665630500165,-0.00332185972365229,-0.0078778935350593,0.00737934665144002,-0.0150917261893305
"2194",0.00516765085037219,-0.00219263747697684,0.00608167852039587,-0.00177348275588685,-0.0162979373484763,-0.00569096261844104,0.00874841581637775,0.0043827934431897,-0.0062265360885132,0.0113257646300211
"2195",-0.0129798627887578,-0.0302732212309329,-0.0146804386689416,-0.0186557210214856,0.0139038424801206,0.00497300200352102,-0.0132155130635744,-0.0148871179264426,-0.00681837286297216,-0.0059289081563676
"2196",-0.00159886340760063,-0.00377658033853157,0,-0.0159926245091431,-0.0000818325119624763,-0.00112022865897254,0.00460380998620646,-0.00338714468094781,0.00398923829678788,-0.00795224601006539
"2197",-0.00361586903246436,-0.00404317130477838,-0.00701147604992203,-0.00429317914491001,0.00681615637686561,0.00149523155570108,-0.00916549045117376,0.00967301503252793,0.0209757621421571,0.00601201054571754
"2198",-0.000258842562503525,0.00659710919100509,0.0247132415039764,-0.00215587919062543,-0.00864613728894215,-0.00261312608339481,0.00503662770639779,0.0137238298254974,-0.00615440322480598,0.00597601393501157
"2199",-0.0250973690687439,-0.0186537512087048,-0.0241172266571912,-0.0212964531140641,0.0171137149527718,0.00570784962980508,-0.0180181605778001,-0.0153260320692158,-0.0126582280786489,-0.0138613336739144
"2200",0.000585045492378589,0.00436661332499977,-0.0123565016986178,0.00473049436454565,0.00283121367893124,0.00344254745419303,0.00702428891169116,0.00337244542355908,-0.00405824578598513,0.00669341801839107
"2201",0.0186584477395648,0.0179028088553228,0.021447877400584,0.0288762107932132,-0.00346839045396774,0.000185540312183319,0.00996409468788007,0.0170631765806379,-0.010372309398806,0.00731379861976911
"2202",0.00260933007789421,0.000251584616074441,0.00699892326073082,0.0054913122237441,0.00426620843727155,0.000779676110946648,0.00465109367347094,0.00152492920090075,-0.00121652628470403,-0.00660057038275963
"2203",0.0149377562550621,0.0198438189875771,0.0121632632875579,0.0266988029233171,0.00605794845251584,0.0048242466730759,0.00869852629604306,0.0114212117306238,0.0211748799444895,0.00664442739342297
"2204",0.0177948492279514,0.0189657321351868,0.024892794561189,0.0215722965557883,-0.0135676576372561,-0.00553958560174594,0.017941331880136,0.0225848744451178,-0.00201854302263582,0.0132014125057576
"2205",-0.00342604107737932,0.00459278912865391,-0.00837517838415092,-0.00173564826746997,0.00431329989009144,0.00204257704774347,-0.00245945958661609,-0.00319002192997919,0.0100211825876946,0.0195439748149826
"2206",0.00819018503758762,0.00962449083946959,0.0160472556337674,0.026659051779975,-0.00332255707656515,-0.00250178713529992,0.00972473486368486,0,-0.0014564354500598,-0.00191690668555067
"2207",0.00902676699108285,0.00881808348021385,0.00332495917271536,0.0107253553344606,-0.00837434504339263,-0.00260104195191702,0.00827469606991627,0.00960094932497157,-0.00510481326631207,0.00448137263945814
"2208",0.000596198264691594,0.000944933704173589,0.00248555033317666,0.00363028584191949,0.00262370443383908,0.000559213943311709,-0.0010762363078326,-0.00414518859457313,0.015851237088613,0.00446151072916767
"2209",0.00094375774932165,-0.00354026975672717,0.0016528731041372,-0.00751286061466849,0.00760527851543169,0.00335076669205336,0.00538697920176934,-0.00195912563289902,0.00396856668254975,-0.0158629878376184
"2210",-0.00630187558265216,-0.0106583556531175,-0.0107260021949709,-0.0162598926227694,0.00170437460980732,0.00092725734577126,-0.0073675430645308,-0.00981325524367049,0.00494118237249452,-0.00644743147882887
"2211",-0.00479418855958313,0.00526687958461358,-0.0116763939386997,0.00769453199000036,0.00875054444946577,0.005468388710542,-0.00647778053280712,0.0094150892502225,0.01743247794178,0.00259568152702783
"2212",0.0153544235553931,0.0126218523402915,0.0253163384090249,0.0243212107839732,-0.00489935645876549,-0.00341053519918522,0.0114100918799778,0.0130093894712688,-0.00456899226024055,-0.00258896140772769
"2213",0.00454668170826422,-0.00188147621264889,0.00493845800636539,0.000828244501405617,0.00032281795900202,-0.000832463598635869,0.00805786971894884,0.00315004926578366,-0.00706154994208186,0.000648920381757012
"2214",0.000492017556591895,-0.00376983223344773,-0.00491418948794387,-0.0102067559420689,-0.00274352641026787,-0.00046287407747525,0.0118570389665424,0.000966202342952416,-0.004178158132779,-0.0181582545830651
"2215",-0.00127839813621911,-0.00307471324471931,-0.00576121608773472,-0.000279017339173238,-0.00614927001997234,-0.00342664409661131,0.00118522888808803,-0.0012065241142265,0.0063382076326961,0.00198147886929001
"2216",-0.00620371909440498,-0.0045078781082698,0.0132450999617693,-0.014496641046729,0.00993227020846388,0.00343842635999936,-0.00355111943143738,-0.00507366139031873,-0.00887075289086969,-0.00856956398348829
"2217",0.0168938921451018,0.0102478613577182,0.0122547233144297,0.0206507240412339,0.00169276153267339,0.00101881071931986,0.0109543800091279,0.0179696651615384,-0.000358014847632204,0.00332449124458023
"2218",0.010961488619877,0.00825666184375184,0.00968533441098152,0.00582039252104161,-0.00853043590114211,-0.00564355102740344,-0.00913840084372952,0.00238563626662924,-0.0017011549520789,-0.00596420155884292
"2219",-0.00245750886118767,-0.00491359814382897,-0.000799254032444963,-0.00909357435704283,0.00665591120313658,0.00260478849305934,-0.000131551920563688,-0.0038079709644,-0.000627802690582935,-0.00266663025528879
"2220",-0.00193243236451057,-0.00940477088083047,-0.008000055767866,-0.0114014830781868,0.0024995229756557,0.00250595794984831,-0.0025036510928752,-0.000955460227845317,0.00224356097998735,-0.00467914912177814
"2221",0.0113746396683967,0.00735792700218063,0.00967736987739065,-0.0115331010191829,-0.00402137560976512,-0.00518365006731869,0.00383085237141345,0,-0.00805874820916908,0.0167897693851011
"2222",-0.000574349334119262,-0.00424116798418439,-0.0111822136101104,-0.00939085819740304,-0.0159087594309425,-0.0061416994674458,-0.00105272599412876,-0.00645624253340094,-0.00956849620480682,-0.00594450458779516
"2223",-0.00430975759834784,-0.000709961330592424,-0.00484644815128099,0.00172361788628517,0.00754939551150158,0.00196668202777706,-0.00724543789538701,-0.00216613880236383,-0.00382790736576821,0.00996670947658385
"2224",0.0118311285615784,0.0113663792181171,0.00730516348776766,0.0197876428670234,-0.00459524182632021,-0.0028731829077574,0.0221601925382298,0.00554762467954251,-0.00649594675674436,-0.00526308626300498
"2225",0.00289915114061001,-0.00210723110898059,-0.000805694481556984,0.0132171235855298,-0.00820034573535267,-0.00262764428149687,-0.00986641089216445,-0.00407779615879245,-0.0148263473552389,0.0178571708144006
"2226",-0.00303310395472567,-0.006804201831349,-0.00483880459692088,-0.008048851842135,0.00115756346999452,-0.00103557623396289,-0.00432648374746458,-0.0144505217255252,-0.00944103544285746,-0.0168941229624917
"2227",-0.000998315784505044,-0.00307094760198834,0.00729332381586012,0.00167876740509398,-0.00264256629820736,-0.000659093515096409,0.0028970582660075,0.00171049647723365,-0.00311410773696219,-0.0079312219733344
"2228",-0.000523492275505966,-0.00545048814594695,-0.00241338970956828,-0.0139664166095658,-0.0146559431637032,-0.00678659393698844,-0.0286239908790491,-0.0124419822706928,-0.0145778210391692,-0.0059960575746596
"2229",-0.00933157073559943,-0.010483752890379,-0.00403228640000508,-0.0249291585143203,-0.00563019920467478,-0.00170845626839267,-0.0135172876920917,-0.024950591929327,0.00288188286036273,-0.00871308670317672
"2230",0.00230692959976597,-0.00433412696309399,0.010526333264772,-0.00435788534289416,0.00295773400868415,0.00190159329806239,0.00918078912833864,0,-0.00210729881020499,-0.00202843934733932
"2231",-0.00393160574664819,0.00507866115338063,0.00400643845496096,0.00204270857604927,-0.00210684034713604,-0.000474780437188516,0.00122180802813321,0.00810748100571446,-0.00335955077750061,-0.0101626021929274
"2232",-0.0139600340553065,-0.0153995994720076,-0.00957713827991991,-0.00961008227173354,0.00481334998783867,0.000569578781451474,-0.0071873473570675,-0.00804227838645355,0.000192584027880471,-0.0143737315317003
"2233",-0.0112282124465952,-0.00855327246426307,-0.00483473209066154,-0.0138192641785628,0.0057142244863746,0.00379504064885117,-0.0105176766113503,-0.00481407421948576,-0.00279248922084718,-0.00763885608064085
"2234",0.0152069523144807,0.0125708810217,0.00971663716545068,0.0193797933889139,-0.000918896307229744,0.00132360973973777,0.0117337245996016,0.0132385824741643,0.00144844537366651,0.00489846340708389
"2235",-0.00072954897176214,0.00316472304187387,0.00240582102855802,-0.0029246818209181,0.00167250357041859,-0.00028352103556939,0.000546061016041932,0.00477383052862268,-0.0132099413095164,-0.0153202689780357
"2236",0.0158660113794353,0.0101917185122535,0.00480000756232979,0.0108534064266399,0.00208737813481297,-0.000471976113383676,0.0106365611054218,0.00725182299435367,0.000879460655831998,0.00424322340568328
"2237",-0.000862235583119042,0.00576498979080142,0,0.00899620136762369,0.00666548836566627,0.0021727475014155,0.00283373883062232,0.00570975153142816,0.0110319047154153,0
"2238",0.00364411338274495,-0.00740380760371384,0.00477692720169642,0.0100659659796767,-0.00306244434249825,-0.00131975504271342,0.0102259395793893,0.00444362803153719,-0.00453845122708474,-0.00140843151233594
"2239",-0.00114649309122483,-0.00697804397786905,-0.00475421665483533,-0.00939639485606936,0.00307185171741109,0.00132149909781165,0.00173176868573433,-0.0105677193382328,-0.00805115949369128,0.0077574441065984
"2240",0.00133903903820776,-0.00169605908871551,0.00477692720169642,0.00517392250393045,-0.0000827687660135412,0.000942412114327107,-0.00491946963700618,-0.000745333067086573,0.00664971627909816,0.0160951672652541
"2241",-0.000143053022727768,0.00582526897442115,-0.00633906954925956,-0.00772074575908976,0.00231759745190474,0.000565009317634591,0.00333988402909458,0.000248737838009605,-0.00466293948585716,-0.00137739162486072
"2242",0.00114643291536565,0.00482622180509673,-0.00478469681817928,-0.0219021702635001,-0.000990780731721985,0.00103530993458878,0.0079905677888723,-0.00472150204057054,-0.0118094769842814,-0.0151724188841127
"2243",-0.00415166795727717,0,-0.00801296337623991,0.00147319419476455,0.00396760574187116,0.0003759136904955,-0.00634132955990718,0.000499254996543019,0.00661726419753084,-0.00630257884926444
"2244",0.00953584582313138,0.00696452947990722,0.0153474489989149,0.00764937350870309,0.013507564064412,0.00531843686535516,0.0123652108177357,0.0187171835061164,0.00353219198454058,0.0112756100009341
"2245",-0.0102051013978794,-0.0114477017006201,-0.00795539841506265,-0.0119710146468306,0.000325719107506339,-0.00280883520054898,-0.0189127006885078,-0.0142087092120182,-0.015545532025279,-0.0209059238447552
"2246",-0.0140027294505882,-0.00506619019628884,-0.0096231326768349,-0.00561445207104205,-0.0271833581316751,-0.0105163833459285,-0.0147256673593718,-0.00670983928296709,0.0106266757249642,0.0113878176129558
"2247",0.0195028689356465,0.00994161382070557,0.00566785085112587,0.00683496331493938,0.00878451863069118,0.00370092646054809,0.0167121531951315,0.00850644766699227,0.0222090699251363,-0.0014074403706511
"2248",-0.0060585191319491,-0.00672266513327857,-0.00241541990233729,-0.0165288649611878,0.0097032109702988,0.00321471255712669,-0.00267291352745447,-0.00868261863414865,-0.0129782641697249,-0.0288936282311872
"2249",-0.00671953484113941,-0.0157117065966428,-0.0129135542207369,-0.0111044217583951,0.000492606840332144,0.000565265951348204,-0.00241152874752937,-0.0102605240433068,0.00165577094878278,-0.00507975678233286
"2250",-0.00777967337888075,-0.00221043425296319,-0.0114471699849166,-0.0081941668466905,-0.00106726217589226,0.00150691037891648,-0.00617873355074805,-0.00278137704983838,-0.00194473947665263,0.000729459707354385
"2251",0.00258111889293722,-0.00319955110916903,0.00909828687358782,-0.00673210969364346,0.00131511702102194,-0.00216314630597403,-0.00567642876688423,-0.00329584685031947,-0.000876812167544982,-0.00364433985582713
"2252",-0.0193811009477631,-0.0170368201626206,-0.0155737092468744,-0.0280345212523885,0.015758406110814,0.00801162718933823,-0.00462128738172007,-0.0167897473324921,0.00546073119081236,-0.0102415653600367
"2253",0.00505242233924474,-0.00150719389991216,0.00915898218077094,0.0161648871408626,-0.0129285050326116,-0.00738697223347617,0.0031404874438028,0.00491587289609607,-0.0128018619648738,-0.00665179463204035
"2254",0.0104980891382007,0.0090563579992069,-0.00412544196235187,0.0152838034807081,-0.00589400913551685,-0.00254326344928713,0.0110261334385051,0.00334736564572347,-0.00265255916443108,-0.00223211243083221
"2255",0.0146319284220169,0.0184494333269769,0.0248551010161888,0.0196622104050981,-0.00214074443702195,-0.00264416687869862,0.0196584631346122,0.0207848492710911,0.0121158691523602,-0.00447421180545382
"2256",-0.0152383913765709,-0.014198321074159,-0.00970092734747641,-0.012955930090176,0.0113055164663722,0.00416623249626924,-0.00488581559997781,-0.0145799192816276,-0.0218978102189781,-0.0104869787599111
"2257",-0.0178148677972114,-0.0124162175809316,-0.0122448969704209,-0.0033575307149285,0.00554857944485754,0.00358319690875564,-0.0127389789201766,-0.00282342810557523,0.015323393034826,0.00454210752137274
"2258",0.00824892011672085,0.00475441551094047,0.00316363501699124,0.00780741925835304,-0.000243133456957256,0.000470107449640045,0.00510734520857392,0.00360361943008103,0.0108780967181683,-0.00452157006397669
"2259",0.00907448873558603,0.0072992388403792,0.00746886830648608,0.00802459516454834,-0.00722400679005397,-0.00281766359712277,0.00414545542814149,0.00487288741932557,-0.00523510411565486,-0.0045420296094798
"2260",0.0123831414436784,0.0194902312538829,0.0107083907105192,0.0140844528320503,-0.00752230725930847,-0.00226011688081917,0.0113201220540826,0.00995420975422401,-0.00292372085641046,0.0182510150888562
"2261",-0.00165030726865067,0.00147060771321961,-0.0122251242683519,-0.00362315312971428,0.00572934253455037,0.00183363429413252,0.000266408878899949,0.0015161616576298,0.0072329685706769,0
"2262",-0.00228511022473676,-0.00416045169626511,0.000825159992828173,-0.00696953777337306,0.00295512967337852,0.000188761733996401,0.00293372072413134,-0.00656055698025071,-0.00756919919740318,-0.0141898071176862
"2263",0.0106719766013514,0.0088471944516828,0.0148392430242072,0.000915337288331264,-0.0166138695841486,-0.00528320337008292,0.0102363251638173,0.0104139041183904,-0.000684462716861178,0.0166667524346811
"2264",-0.00708779981647967,-0.00803874107681501,-0.00568648873967359,-0.015548803104815,-0.000998339945373572,0.000379312679735122,-0.00447415343827873,-0.00703864678456201,-0.00763208437276164,-0.00968705542198245
"2265",-0.0100032776368154,-0.0149805357157816,-0.00980394495034864,-0.00309702224658992,0.00449829413849101,0.00113790836142758,-0.00753486871204367,-0.0096204694989096,0.000394409394486317,0.00526712378627625
"2266",-0.013979536148481,-0.0149589773104761,-0.015676448895698,-0.0273375535366791,0.00721524035306542,0.00426136721763437,-0.00972281009925713,-0.00894695485623631,0.0140942244637712,-0.00748492787745059
"2267",0.0016912689914137,-0.00632735446862465,0.0125733339909304,0.00223579895328263,-0.00403457953282871,-0.000282766119730993,0.0164092310522321,0.00154815034036115,0.00281855382270924,-0.0098039421145949
"2268",-0.0126142208531249,-0.0168111397738384,-0.0173841182014508,-0.0191205480743303,0.0134753944674944,0.00603731641525185,-0.00330850957809936,-0.0100438301498822,0.0144407637138981,-0.0159939228439159
"2269",-0.0239915768024475,-0.0181346656092086,-0.015164280894201,-0.0308642939863112,0.00179483858307194,0.00215641421206691,-0.0223050507448107,-0.0228929756493788,0.0141397155658682,-0.00464405853976857
"2270",-0.0109764124444166,-0.0100263404236193,-0.0213858817272133,-0.0107274612447024,0.00447825364397159,0.00252633735951302,-0.0118139066910531,-0.013578347272067,-0.0044277154135145,-0.00466564641415823
"2271",0.000989880026305068,0.00346493973090278,0.00699321883096804,-0.00033885562809266,-0.010943749559469,-0.00317341708134888,0.00398513350978358,0.00377869448642731,-0.00889479560938689,-0.027343700059397
"2272",0.00806845318544247,0.00796802289133547,-0.00520851907234643,0.00203389704901502,0.0144254863586135,0.00449420603867301,-0.00698069584609895,0.00430228099671792,-0.00506013948940498,-0.00642569783124736
"2273",-0.0249407691781877,-0.0171276854501491,-0.00872605145266192,-0.0104871999582878,0.00985673308793267,0.00391460833190505,-0.0151620408990426,-0.0109775019502681,0.00489398334990865,-0.00565877484512667
"2274",0.0164168550263235,0.0128684998380684,0.0123240638616968,0.0129916076488972,-0.00936048535023226,-0.00204230115485149,-0.00139934268372743,0.00893357548008433,-0.0162338042758421,0.00243899091980437
"2275",-0.0214660752997756,-0.0367920092116133,-0.0278260423244094,-0.0394870889233299,0.0155869721984294,0.00465133967071862,-0.0113524814802886,-0.0300508370576997,0.0102893130544353,-0.0210869089061161
"2276",0.00133123320812034,0.00906849976457935,0.00805007766095378,0.0147574683883072,-0.0031014421953125,-0.00129620329013991,0.00297724735277027,0.00553247645153121,-0.000960789758632008,-0.00828489181420122
"2277",-0.0128151192954098,-0.0206971352927823,-0.0381544767233861,-0.0218142790489818,0.0105296411832807,0.00491398543231147,-0.0265729084319444,-0.0220081819502859,0.0133679549903456,-0.0075187801837816
"2278",0.00560204487021876,0.0108454800856879,-0.00369001265020841,0.00389389298329634,-0.00678886512426657,-0.00249114176100884,0.00667941388578286,0.00450053506539771,0.0011387965890064,0.0134680023834841
"2279",0.0205151317742818,0.0264097236004661,0.045370486459378,0.0342030641873465,-0.00381497023319544,-0.00221969958252488,0.0276935680192065,0.0229629005747729,-0.00464497117537155,0.0299002652026497
"2280",-0.0151166718804302,-0.0134011998189386,-0.0212578685755503,-0.0170474664264765,0.00542539901182626,0.00333699670719434,-0.00982430421468183,-0.00848627622642451,0.0102857333333333,-0.021774146157322
"2281",0.0136433033074772,0.0214614921821286,0.0135747711780834,0.0145680729481956,0.000476327774119767,0.000739149841444187,0.0214031063657585,0.0168415148217682,0.0114064760292898,0.0197856396611851
"2282",-0.010883361135584,-0.00851066186933813,0.000892821275057187,-0.00341867693316134,-0.000238222006286648,0.000738463451070315,-0.0155424250452442,-0.00705949903077385,0.00372822253958227,0.0121261125018888
"2283",0.00520922952583591,0.00214619298378405,0.00178407360311206,0.015780460119674,0.00142809787473097,0.001291730844446,-0.00662580153209091,0.00710968987958793,-0.0106788093475939,0.0111821204449172
"2284",0.0243774244564392,0.016059835732168,0.0240427565844004,0.0324214934055871,0.00847645169806865,0.00534441675617803,0.0217118341726072,0.0285095830663056,0.00384828229915257,0.00947862482423667
"2285",-0.000361334735548557,-0.00158072100487816,-0.00608685215063798,-0.00948639397707429,-0.00306141471088861,-0.00230391189893953,0.00013870950022965,0.00712780477204733,0.0102852363801376,-0.0187792482003014
"2286",-0.0180224132214298,-0.0274404043199921,-0.0104986872950545,-0.0323646210806806,0.0185522480810896,0.00708364031580166,-0.0105541699779617,-0.0212321442436937,0.000370134186854276,-0.0175439474833902
"2287",0.00599522956648935,0.0151927582462399,-0.0123783783732585,0.0283276370550229,-0.00829336430228189,-0.00109623860506491,0.0049122996888491,0.0182108409046635,0.010731834979437,0.0251624127265246
"2288",0.00156805843957741,0.00133591532674249,-0.00268604094276359,0.0076336307121172,0.004845589073047,0.00237778200117078,0.00111758894638303,0.00236733473935069,0.0120823798627001,-0.00158359108553852
"2289",-0.0190500110064732,-0.0152120250867369,-0.0170554542308498,-0.0115284740484218,0.00116665730759369,0.0012773031896538,-0.0224612166779103,-0.0170561488495028,0.0158270778692231,-0.00634416643820135
"2290",-0.0134610796627123,-0.023577436866375,-0.00182650845372834,-0.0136620800523344,0.0215195863085742,0.00747166226403539,-0.0293989080003992,-0.0149488991447826,0.01344375,-0.00478852442938482
"2291",0.000054061447636089,-0.00888154296209476,-0.0192131872350615,-0.0138512809369771,0.00106464664387995,0.000180645060755991,-0.0161741255598917,-0.00406516114805977,-0.00219625753850028,-0.0256615684840983
"2292",-0.000862995058011573,0.00420060730190452,-0.0177238685485288,0.00411099399176229,0.00881284955425388,0.00298400507115826,0.0052309959893404,0.000271860381546585,0.00774781638056332,0.0016460680853132
"2293",-0.0130079227837007,-0.0142218954632493,-0.0199431346465897,-0.0167178567560625,0.00700342750217309,0.00459803335191378,-0.0147192876790483,-0.00843272306558784,0.0401887038283129,0.0123253916243458
"2294",0.0206168453482016,0.0195191760306186,0.00872104814303509,0.0173490258013167,-0.0166019513474404,-0.00762808972507401,0.0129772399014374,0.0150893021588874,-0.00587936344497497,0.0146104412805887
"2295",0.0168781077222806,0.01609287759583,0.0365033111683206,0.0221691283476813,-0.0105701408360324,-0.00298442164691948,0.0192165351559719,0.0202703776067124,-0.0303312265095367,-0.0112000939303752
"2296",0.0163347622186762,0.0207540261821471,0.00834097017973834,0.0196863164980472,-0.00614885083717631,-0.00244900044746654,0.0090616207732761,0.0127148564539392,0.00618633805488367,0.0210357295389787
"2297",-0.00409580935022813,-0.005885727790782,0,-0.00589001314610849,0.0122962635879056,0.00463725402567139,0.0095597173918065,-0.00392373704279092,0.0243331999220679,-0.00554667519181595
"2298",-0.000468503326832792,-0.00188369527600141,-0.00459562583676154,-0.00460830405041557,0.000839921924084441,0,0.00215216739202639,0.00787821643664732,-0.00600218948345443,-0.00876506550734024
"2299",0.014479312180814,0.00727976252123419,0.0166206995279345,0.0248016443555237,-0.000533893605510039,-0.000995617669813154,0.0115962038368289,0.010422281810573,-0.0177751655421812,0.015273351601643
"2300",-0.0126296056627673,-0.017398499411745,-0.0163489682392385,-0.0212971783698916,0.00404734162257903,0.0019932198245034,-0.00240582258670574,-0.0167613014152151,0.0149796781536007,-0.0134600760332335
"2301",0.00457559287687337,-0.00435832869427955,0.0101571092680075,-0.00230796837442904,-0.00197777610861205,0,0.000425456975914118,0.00550731151470241,0.00332707726218162,0.0128411642829631
"2302",0.0121118721685456,0.0139534098620515,0.0118828885929345,0.00330478680411628,0.00358240270224019,0.00298396068524442,0.0181511306023727,0.00834626759679424,0.00263580475609393,-0.000792463724620274
"2303",-0.00230150879215041,-0.00296803188275385,-0.000903233641757706,-0.0098815234669124,-0.00964470050206989,-0.00486812137890125,-0.00306429109322026,-0.00646633394639218,-0.00686903844757536,-0.00158593958574915
"2304",-0.00784244964585445,-0.00460107016341793,-0.0153707423103369,0.00864941075439241,0.00437091829963543,0.00163069772620528,-0.0016764191320412,-0.00104149171096768,0.0130646228924549,0.012708406021543
"2305",0.0235068700351397,0.0274607439212458,0.0247934028600945,0.03562002794313,-0.0176087788856392,-0.00781626223771181,0.0260286129205112,0.0242377045696183,-0.00733312548325293,0.00078430302575816
"2306",0.00449262984725451,0.00238177767880354,0.0143369185948776,0.0133758567998801,0.00412689640004849,-0.001734587595556,0.00763765607405276,0.00585235607680978,0.00772695103320764,0.00548589929572096
"2307",0.00391956776358948,0.00844751246289599,0.0070670673356219,0.0113135622245235,0.00364447131171497,0.00118899169113651,0.00500818487919363,0.00455371176103814,0.0172733653522075,0.00545596840250417
"2308",0.00325360475335268,0.00523570069372581,0.0105265052121097,0.0198881728255198,-0.00641266697356158,-0.0033793440341936,0.00269364863885024,0.00302192650534883,-0.00157377615570831,0.0193798199127144
"2309",0.000798322477178592,0,-0.0104168521635167,-0.0015233381174814,-0.000311186472022662,-0.00201609285894477,0.00188017794751461,-0.00577464332663757,0.00497758416311944,0.0182510150888562
"2310",-0.0109177725879248,-0.0106770913271598,-0.00964897146673926,-0.0170889645734349,0.0110457163558544,0.00578489423903061,-0.0103229115630816,-0.00303035376724592,-0.00462272580999457,-0.0134429144816003
"2311",0.00493932484360382,0.00552767996254167,-0.000885893770173674,0.00620929295989736,-0.00607824333917029,-0.00392555257334393,0.00406380305162779,0.000253390178182489,-0.00829324915751783,0.0151400727276354
"2312",0.000802444987857642,-0.00052356712218915,-0.00443256538921322,0.00154267643704076,-0.00410216591719836,-0.00357469983068104,-0.0025633161520302,0.00177265763571022,0.0160561796946617,-0.00149140393515124
"2313",0.0161372447988211,0.0267155274696498,0.0267141845817738,0.0209488579569388,-0.0101042795139561,-0.00285154126298603,0.0236710824255626,0.0245194962492099,-0.0172016131687243,0.00373407885778065
"2314",-0.00128226398411513,-0.00280611652181595,0.00433645562629081,-0.00603510911617133,0.00314078340353885,0.000737927655383386,-0.00132129846926254,-0.00197361302215149,-0.0128967502588812,-0.00892852630190855
"2315",-0.00162966417705035,-0.00946530326270378,-0.0129532190467452,-0.0142681711065537,0.000939092105588291,-0.000184782842755804,-0.000264649513843196,-0.00296696346565961,0.000763519111813382,-0.00825829985097226
"2316",0.00578699765622193,0.010330511349161,0.00174973435444326,0.0200183742214184,0.00297154730433191,0.00525605105332438,0.0127051478107034,0.0126457107213724,0.0222956682120692,0.0174110485764289
"2317",0.00634424479312812,0.00741314311587216,0.00349333287364639,0.0220411699953849,0.00413243523768947,0.00110016254004686,0.0139830162149042,0.0173849303154043,-0.00381457015721265,0.0111607918898995
"2318",0.00392964238340987,-0.000253674639992152,-0.00348117198112596,0.00531754136345408,0.00209632249851666,0.00174070623173961,-0.00386640905965474,-0.001666878183051,-0.00274697417997938,-0.000735900819623936
"2319",0.00141881231467589,-0.00482235554949773,0.00436675380370932,0.00205696426162327,-0.00767081274956904,-0.00283472532026829,-0.00646895142158221,-0.00121003368287842,-0.00701171935696865,0.00294554370651778
"2320",-0.00053755536440947,-0.00535580402611435,0.00608701516720078,-0.00234592198952699,-0.000234357863379109,-0.00210972638189466,0.000260479364800448,-0.000726793302264772,0.00294215705230449,0.00734219461659547
"2321",-0.00659945788914895,-0.00820514984818832,-0.0129646446915489,-0.0170488352310828,0.0113248499983272,0.00459525885933787,-0.00704843666682009,-0.0106694461205585,-0.0226300984432167,-0.0211371111512028
"2322",-0.000442707414448296,-0.00723877505686166,-0.00612958604727454,-0.0023923536471846,0.000386102622693674,-0.00100608913207823,0.000796385137287414,-0.00661791707246984,-0.00240115768457971,-0.0059567318472874
"2323",0.000590669382952491,0.00416648672540698,0.0149781045824349,0.00329730512232085,0.00131260214036111,0.00146519730708516,0.00768909516113592,0.00320758984179026,0.00232094898442448,0.00299621356440394
"2324",0.00925006118629379,0.0121887104306468,0.0104165034488115,0.0137435983588492,0.0104847352095392,0.00676732163963156,0.019865420763356,0.0150027140339011,0.0185249059781287,-0.00224052417919829
"2325",0.00438773410210125,0.0107610392935442,-0.00343631147224333,0.010315488432237,-0.0105290581547435,-0.0013625775712115,-0.00154768694505003,0.0082382225943618,-0.0139778037390064,-0.00374246393872524
"2326",-0.0024269361765763,-0.00861853331399198,-0.0163794834997236,-0.000875145206503336,0.00709401766626416,0.00363850778065,0.00594309768917523,-0.00360501918914258,0.00461145182940137,-0.00150268636214512
"2327",0.0068120398103666,-0.00869325667020604,-0.024539764261697,-0.00291972713170574,0.00260840071181656,-0.00029089850028452,0.00064239320950632,-0.00892409039597541,-0.00603535367252084,-0.0173061642997535
"2328",-0.00323795930421777,0.00128951418532397,0,-0.0120059224915666,0.000612095000930291,0.00118049284343535,-0.00141216511835218,-0.00292041216299888,-0.00667064055417776,-0.0137825107354482
"2329",-0.00998798104363585,-0.0190621861805117,-0.0215633676774732,-0.0195613386255007,0.0109359595353875,0.00399028919847377,-0.0056554168371713,-0.00610182311441976,0.0130004474730874,-0.00232932034986943
"2330",0.0109212262466767,0.0152309967243491,0.0165288532648782,0.012091912332892,-0.00726214726965246,-0.00216788782724664,0.0024560208629314,0.0098229368287206,-0.00611934366413924,0.0108950335716682
"2331",-0.0119656894454048,-0.0168132475420067,-0.00541988570411089,-0.0200119881257546,0.0123449838188083,0.00515979608183637,-0.0054156932200472,-0.00851165469150916,0.0142808189792916,-0.00307932878634831
"2332",0.00269652213076044,0.0176269512506628,0.0290642675560357,0.017372774335672,-0.00632292927215572,-0.00153105004068754,0.00570454193844494,0.0129995994777803,-0.00151758703720095,0.0239382940858939
"2333",-0.0023471309782831,0.0018097883590491,-0.00617808805420639,0.0128819130084703,-0.00128798542545783,-0.000180153500774383,-0.00128924723125989,0.00411630827247067,0.0135100819049228,0.00754137452184356
"2334",0.00931277622733484,0.0113546974533281,0.0230906337145482,0.0153802064975663,-0.00690247008005218,-0.00396963444452147,0.00684169551409397,0.00795757398371189,0.000166658336804515,0.02170659899314
"2335",0.0101012362518995,0.0137791221530676,0.0277776602480067,0.0177686914057749,0.00351386234778528,0.000724821518029106,-0.00230779786019475,0.00885181035962423,-0.0106622737860324,0.00512828594201653
"2336",0.0000479453667721064,0.00125846893543202,0.00422300718853785,-0.00486539670820263,-0.00479530244114545,-0.00235334933858145,-0.00642525939232408,-0.00545437777414004,-0.0139765600903401,-0.0080175326796712
"2337",-0.00110594156149357,-0.00175965903549635,-0.00925150592395863,-0.00575218522206178,0.00856531890546464,0.002993928144017,0.00659623105107054,-0.00238423056112946,0.00691654848504375,-0.00367379462428574
"2338",0.00702685597260189,0.00906576110836199,0.00764005706552329,0.00462827656814868,-0.00432167381238946,-0.000995124301886641,0.00423973699798696,0.00693127513906688,-0.0015264586419006,0.00442479420991582
"2339",0.00315431882792594,0.0197154342883619,0.0151643937050379,0.01526058139409,-0.00312244303852371,-0.00162965289300365,0.00102355902270612,0.00593384708468081,0.0156276883918411,0.0212922283683834
"2340",0.000952830638455859,-0.00244730345711486,0.00580891729824384,-0.00453773727451678,-0.0110005960412526,-0.00507836705441367,-0.0140593022967882,0.00259565005525864,-0.00510119576683066,0.0194104523215852
"2341",-0.00537843924345516,-0.00711478769793683,0,-0.0099714512359006,-0.00594828060661856,-0.00164071381804187,-0.0169821209707509,-0.0112967513140242,0.00378244091970714,-0.0042313265506686
"2342",0,-0.00222385697434735,0.0074258433224399,-0.00604325533661298,-0.00256412841774234,-0.00109535986632503,0.0106816174616151,-0.000713929529663537,-0.0128119161415494,-0.00424916097384553
"2343",-0.00172279023040067,-0.00421010194171156,-0.00655202898889595,-0.00636944368385661,-0.00412900161154839,-0.00109708504580464,0.00626327704366458,0.00905181566639612,0.00288407840261318,-0.000711300967053075
"2344",0.0014861254373788,0.00547123603579913,-0.00412197883332865,0.0107808045966029,-0.00453755017723012,-0.00210422592982873,0.0036306626700453,0.00779047273012634,0.00397525152731326,0.0128112856578488
"2345",0.00205810863079559,0.00469950103966776,-0.000827781369678204,0.00605377193917267,0.00998069254118072,0.00550145223654241,-0.000258230814461746,-0.00163978495356143,0.00286439771350633,0.00913564938547906
"2346",-0.00907590810673597,-0.00516989383495758,-0.0455674466412721,-0.0103152415648027,0.00412367223533838,0.00346537069952491,-0.00232639354911235,-0.00633519099370816,0.0189012095186389,0.00557102644813079
"2347",-0.00539859880522753,-0.00247455633378846,-0.00868069463783261,-0.00434269318500169,0.00255762461297482,-0.000363624287424535,-0.00829008851903079,0.000236218554778178,0.0194575066414584,0.00969530142169384
"2348",0.00794841418719328,0.00744211278874052,0.0183887112393841,-0.0026171650094583,-0.0100683541759813,-0.00290422047988459,0.0133226219301201,0.00873442202945829,-0.00331584305190713,-0.0137173754198485
"2349",-0.00870324438420256,-0.0201917588335341,-0.00945808037617057,-0.028279791297329,0.0125956555017233,0.00593507909398094,-0.00219118682489972,-0.0109992756259568,-0.00227198153638397,-0.015299103572847
"2350",-0.00557804914045512,-0.0130686959677399,-0.00868069463783261,-0.0162017724528839,0.00548573196681645,0.00181520072721386,0.0134350993289967,-0.00567902581027546,-0.00609954461694495,0.000706277775116781
"2351",-0.000195127428708308,-0.00483843422569086,0.00525403475306629,-0.00030482639796614,0.00668478307045772,0.00271798995803119,0.00382400276971495,-0.00023795064209764,-0.00114556092910212,-0.00988003858289233
"2352",0.00365901548923797,0.00307066513994769,0.00522648083623678,0.00152533034763147,-0.00427435387256558,-0.00234913850280272,0.00977794252012609,0.00166611246496018,0.0090931432784469,0.00641481120450282
"2353",0.000826450540746926,-0.00127545529173068,-0.000866609144910213,-0.0127932010388226,0.00314295393458486,0.00190187326430191,0.00804833992843501,0.000713079886509371,-0.0205390323104401,-0.0219545936385844
"2354",0.0124336704748904,0.0102170470806375,0.0251518142722733,0.0191297274525142,0.000076459070313728,-0.000180599087817312,0.00187109126758456,0.0121112645699533,0.00273519266083389,0.0246197266652655
"2355",-0.00935483794280645,-0.00581545787507831,-0.0186124989147007,-0.00242191794204583,0.00565448689339587,0.00153698109502698,-0.0178060380258557,-0.0114970142686147,0.0094230448977588,0.0233216012391908
"2356",0.000290537376831823,-0.00279743818317868,0.00775853988403696,-0.00273134309840006,-0.0045591021787621,-0.00270824324059704,0.00494400045059362,-0.00617154456794078,-0.00786111182784688,0.0013812676985363
"2357",-0.00871413444451297,-0.0102014412384764,-0.0136868900783947,-0.0179549918508574,0.00969399527317805,0.00380154347961326,-0.00807360907772037,-0.0100310586059789,0.00453941054673446,-0.00137936242976755
"2358",0.0098652917737303,0.0123679347004704,0.0138768205965372,0.0120855200304915,-0.00861798370865463,-0.00360684096024666,0.00788513139056568,0.012304111287299,0.000739495528218725,0.0110497861959944
"2359",-0.00933346194898388,-0.00865362915329904,-0.00684350231313391,-0.00459287131670061,0.00167766059677832,-0.00135725008524612,-0.0151419113570652,-0.00166806701580058,0.00344825935677506,0.00751355819875688
"2360",0.000292719037028544,0.00333749729238608,0.000861315018280573,-0.00984313066340958,-0.0142355488936493,-0.00806631094629184,-0.0139654365128276,-0.004058299858965,-0.0173457943270676,-0.00745752564579838
"2361",-0.00346502314074204,-0.00614124385532078,-0.00688454425001572,-0.00931962515444762,0.00432445813871873,0.00100509734778931,-0.0107847130551071,-0.0105468167550883,-0.001915029174272,-0.00273227328300718
"2362",0.00631752629130511,0.008238951358021,0.00693226976798655,0.0100345330832161,0.00076872676771722,0.000638803839440927,0.00801274356481607,0.00436048768880082,-0.00133481268036673,0.00410953283883031
"2363",-0.00136254355785981,-0.00306427699481671,-0.0043027998229852,-0.001862638567383,0.00222836955546546,0.0006382383741943,0.000912099970598268,-0.000241164670734983,-0.0028401637527371,-0.00545702180239194
"2364",0.0129622572009076,0.0197234908169068,0.00777856460197102,0.010264173550073,-0.00444605393713893,-0.00164049068371752,0.0119773757373536,0.0125454588598897,-0.0173410400266136,0
"2365",0.0067829984178438,0.0113034865670776,0.006861202536671,0.0120074494669211,-0.00377389416348151,-0.000456624211283896,0.00154383220134058,0.00309738191021691,-0.00272804767106449,0.0116597902841575
"2366",0.000286683138336574,0.00372578985327121,-0.000851777389248687,0.00669301777274689,0.00517910562647761,0.00310591052256126,0.000642475782504315,0,-0.00341939639033861,-0.000677887099525876
"2367",0.00429936608108816,-0.00247455633378846,-0.0025574421030945,-0.000302161869570439,-0.00146108750404939,-0.00191226509373821,0.00436448882618712,-0.00118789143422005,-0.00823467990676474,0.00407050060119052
"2368",-0.0019024250288936,-0.00843477060644759,0.00769222704911066,0.00120914497173041,0.00238737935975908,0.00118607044054775,0.000127780849364934,-0.00784744669362647,0.00380552662673783,-0.00608106773660633
"2369",0.00204908490595734,-0.00125091260201982,-0.000848233218477268,-0.000603809348856621,0.00405726900610293,-0.000337833108495222,0.000639073454449468,0.00143800091446922,-0.00103391351083759,0.0101970756409457
"2370",0.00304370798880438,0.00300616476137194,-0.00848894219078444,0.00815699505868439,0.00720751689394894,0.00310411818159229,0.00536370029156208,-0.0009572700677144,-0.00232882521426903,0.00201895364593252
"2371",-0.00298727017404643,0.00549438081973874,0.00428083357871412,0.0152832779186429,0.0142354342417277,0.00928351771303526,0.0030489507683289,0.0162907944903734,0.0277513534667821,0.00671589392978178
"2372",0.00508867569294869,0.00322901228006756,0.0102301108841361,0.0106257630771114,-0.00743100142002229,-0.00261484079485863,-0.00620565983643862,0.00660089215211568,0.000336482175382402,0.0120079785873621
"2373",0.00156114240195593,0.00693252876816453,0.00675110073940544,0.00905362564034551,0.00242031010015586,0.0014466033513203,0.00611710719938996,0.00491832565226158,-0.00084088464246368,0.00988800541244195
"2374",0.00325983216574,0.00221292091027148,0.00586752742742158,0.00723600182361728,0.00535627306068442,0.00117339532387772,0.00531987688339242,0.00466087741027033,0.0148123379902374,0.0169711811449773
"2375",-0.00136566662116844,-0.0144751519655213,-0.0116667123436496,-0.0114941088173087,0.00645255242952181,0.00153328213217074,0.00151181560257352,-0.00347955323997062,0.00555646034903878,-0.00192551936769392
"2376",-0.00947745888571283,-0.0343538928110562,-0.017706590418109,-0.0252907718399699,0.00484610011932674,0.00351141550693157,-0.00490629242054197,-0.0188547378464026,0.00404122061855672,-0.0122186152959649
"2377",-0.00771180855306974,-0.015210089101762,-0.0180257652605508,-0.0140172981463198,0.00445175144291232,0.00197444116351631,-0.000758597571731578,-0.00972705171784971,0.00739281267279135,0
"2378",-0.00196699287622748,-0.0185863823271325,-0.00437047792040235,-0.00332739140944815,-0.000738682363088383,-0.000269044221417714,-0.00544030747088309,-0.0129372317948746,0.00105999674706458,-0.00651046168649383
"2379",-0.0013939297329808,0.00533458610411208,0.0096575357121107,0.0106222252565686,0.00384424749416135,0.00304566320934496,0.00915909199563525,0.00339798772845712,0.00741225887624641,-0.00524239253493219
"2380",0.00298438824566793,0.00716387433483723,-0.00434776817051308,-0.00360369947819006,0.00485985173879344,0.00107176268324749,0.00504199545235373,-0.000725562734757879,-0.0105110203751617,-0.0171278363614298
"2381",-0.00372410010308466,0.0150156632196461,-0.00174667813171003,0.0027125086425468,-0.00622896158893926,-0.00338979567343733,-0.00150488873793664,0.00383247133077291,0.012828893924552,0.0234584695446547
"2382",0.00643978364611897,0.0254346856002265,0.0227470386524538,0.0177336604622242,-0.0106927596870465,-0.00429643805399404,0.00188448266442576,0.0248055470691819,-0.0059701332626898,0.00916831322138223
"2383",0.00283895493903086,0.0102058203887767,0.00684347940355923,0.00767884428715715,-0.00462092256031299,-0.00224767014537874,0.00411150940065164,0.00783105755119418,-0.0192354761726765,-0.00778717815876662
"2384",-0.00163131963493457,0.00205139537026122,-0.00924826050729399,0.00254016305047422,0.00164725416871092,0.00198240046814058,-0.000503870951716223,-0.00306097663541716,0.000496573998562511,-0.0058862543246091
"2385",0.013022660525873,0.0307061911943531,0.0224719542385388,0.0241601215488481,-0.0114380302290893,-0.00476597309404481,0.00668081330180259,0.0174775540523484,-0.00653433405236836,0.00789483252926959
"2386",-0.0359093158726174,-0.109483705822347,-0.041419977593303,-0.0607017960977838,0.0268468114367069,0.0138235556787212,-0.0121463529698796,-0.0733519253129234,0.0490383727496597,-0.0202349783501855
"2387",-0.0179097556596742,-0.0231391774433878,-0.00529105252705953,-0.0128637641372736,0.0249667286459687,0.00864460839173908,-0.00190121237824437,-0.0230462430585007,0.00539682539682551,-0.00199870871444952
"2388",0.0180361600271361,0.0322488578113547,0.0150707981251978,0.0294756818776525,0.00208400707113765,-0.000176757037573805,0.0217168208979515,0.0358976035796288,-0.0107357120303128,0.0160213488817786
"2389",0.0170275640686621,0.0221179064701433,0.0131006486853331,0.0253166034108148,-0.00767200495569864,-0.00406475798673045,0.0128031856027186,0.0175740799388169,0.00414934567507186,0.014454602712451
"2390",0.0136455676675331,0.0221800393482223,-0.0086208349952257,0.00999407246928352,0.00368460926517189,0.00221833200681898,0.0111682641495057,0.00827046528327169,0.00500639717121421,-0.00582893627845582
"2391",0.00210047767095278,0,-0.00173905372269767,0.0096039923891782,0.013885265668387,0.00264167488754197,-0.00072824829543483,0.000482536498277453,0.0153396298304764,0.0123778149562057
"2392",-0.00719331757885666,-0.0283141997517737,0,-0.021331632949757,0.0125199664754772,0.00548220621711981,0.00765210334894628,-0.0217024025038508,0.00825478519570799,-0.0283139731648793
"2393",0.00599774639244299,-0.00408509899924048,0,-0.0026510535897456,0.00161577469315932,0.000175980759538064,-0.0036158923988675,-0.0014788198201533,0.00587004706982275,0.0039734554960511
"2394",-0.000619884303288853,-0.00519554323595139,0.000870972210665011,-0.00265797223186004,-0.0000701497796582462,-0.00131868585220929,-0.00883144503066868,-0.00271534312658506,-0.00376250491476637,-0.0283641363814513
"2395",0.0148903862070984,0.0156680336541262,0.00696252364129535,0.021616946159615,0.00736628204540857,0.00193672311547122,0.0147684807888888,0.016831907714445,0.0060120161086783,0.0101833702572474
"2396",0.00352700609585455,0.013531988874429,0.0242005784694876,0.00956517657802114,-0.00877509086486572,-0.00527194374614515,0.00721698111130142,0.0131449203027219,-0.00942392707864148,-0.00403234117737061
"2397",0.00726326581148817,0.0149531247608754,0.00590718166245208,0.0140684309651711,-0.0164393308195698,-0.00591891523447652,0.00119386542393451,0.00937044052168479,-0.0165518687900309,0.0188934773809963
"2398",-0.000139602110749149,0.000263106797830481,-0.00167786753442245,-0.00169886693789389,0.0117856309039668,0.00257707059587764,0.00417478828739681,-0.00214237697249842,0.00920176941876893,-0.0125828817108378
"2399",0.00558360700354332,0.0105207224202584,0.00168068750542338,0.0144640663455848,-0.0145428890568049,-0.00416578358511155,-0.00736432724654978,0.00620224437689743,-0.00771512582601408,0.00402422820351811
"2400",-0.00134187082427517,-0.00598662061130439,-0.00335573506884468,-0.00223673022175508,-0.00859625660482533,-0.00382736198354328,0.000837578469497169,-0.0111426552662064,-0.00384831534048036,-0.00267204288248979
"2401",0.00268718813195035,0.00235677197765916,0.00252532019097984,0.00896612671306074,-0.000939457663775012,-0.000268289098562358,0.0025109198473181,0.00311662799342716,0.00157682912572787,-0.00468862042717499
"2402",-0.00101667969767405,-0.00940454906721933,-0.006717105044455,-0.0102749197932618,0.00564115865169956,0.002681406474762,0.00453180718877921,-0.00286786422195717,0.00133814545546174,-0.00605644537272443
"2403",0.00416310138937392,0.00870269836215631,0.00845313962173666,0.00505078031578177,-0.00546597040863694,-0.00205023685632821,-0.000237541662506446,0.0105464524704619,-0.0143070514449103,-0.00677045791683872
"2404",-0.00377709216262545,-0.00235284467865982,-0.00754400793799903,-0.00307119943309142,0.00202481503643792,0.00223310339183946,0.0014250179197286,-0.00189751913205138,0.0152325067009531,-0.00545330161916657
"2405",0.00448515788204262,0.00183427731537855,0.00168920442888099,0.00728079145209581,0.00173221363855358,-0.00080237441700004,0.00830074864038211,-0.000712907230018933,-0.00746272566859252,-0.0020562452815841
"2406",-0.00271601980182301,-0.00026159272880999,-0.00337271165829134,-0.0100081329403624,-0.000720366799375705,-0.000802567215977046,-0.0009408503267887,0.00356720106156239,-0.0069647567386586,-0.0109890024443174
"2407",0.000461382574157732,0.0034015089598014,0.000845986373307017,0.00786289343782021,0.00158608691166817,0.00062467866262117,-0.00459079638453308,0.00545012032145475,0.00422410931518202,-0.00416660978580086
"2408",-0.00106093138858609,0.00651872272929421,0.00169063241664791,0.00334350013311635,0.0124532062120486,0.00428211187794747,-0.0070955700765013,-0.000235756081230609,0.0161111031746033,-0.00976298245846985
"2409",0.00115460384275679,-0.000518027998477111,0,0.000277573548180587,-0.00184849905031348,0.000532724567946508,0.0073842827016195,0.00495068560016376,-0.00288990863774041,-0.00281693550467965
"2410",0.00161454840549924,0.00959049530291134,0.0177215898345422,0.00527502341301633,0.00833405250486963,0.00381787299757796,0.00969518733412156,0.00680268529788641,0.010339902543008,0.00847467913859545
"2411",-0.000828854540970592,-0.0107833181597822,0.00331669126886069,-0.00193312148470437,-0.0108421722506139,-0.00347209004693305,0.00351279493049828,-0.00582482165039011,0.00186079242861803,-0.0175070513551416
"2412",-0.00640756406653609,-0.00259518860705998,-0.0123966526536556,-0.00719428260298793,-0.0103027315037673,-0.00239946071569086,-0.0151691423783599,-0.000937359751211564,0.00812570029309945,-0.0014254239409307
"2413",0.00292293004002775,-0.00416341496780404,-0.00502094348233828,0.00334455287821367,0.000578190905094589,0.000534713194003444,-0.00426530713924744,-0.00821019444653071,-0.00475942259125139,0.0164167665089441
"2414",0.00106387789927287,0.00418082146245857,0.0142977688808279,0.00555548274859063,0.00751394036439179,0.00240401359385234,-0.00238013312363461,0.00709534897707176,0.00169688399677059,0.0042135701416901
"2415",0.00817892818594834,0.00338280686464532,0.00331669126886069,0.0116020827033498,-0.0103976531382658,-0.00621769920221615,0.0013119698655002,0.0023486237935646,-0.0178639569517192,0.00419567454347969
"2416",-0.000595904528366775,0.00103724475521405,0.00413229075220345,0.00710010252797888,0.00188406539156238,-0.000536548717217866,0.000953158770427676,0.00234315071341773,-0.000862414719033699,0.00557102644813079
"2417",0.000596259842306823,0.00958532766417997,0.00905351371033092,0.00677866801818694,0.00983615795302306,0.00357724759065303,0.00368912033993074,-0.00233767319280831,0.00408032793345359,-0.00277004539170966
"2418",-0.00247494166153972,0.00384923998258291,0.00326258532122714,0.000269317577300754,0.00386781109717904,0.00267314952936659,-0.00130420541429965,0.00421743105339822,0.00468895752335863,-0.0118056088131202
"2419",0.00464068302776433,0.00792437671770929,0.00731716084817857,0.0129240551367171,-0.00891827512375842,-0.00479884495667893,-0.00949772694391637,0.000233151597489156,-0.0069228376932613,0.0154603742383221
"2420",-0.000869029223925288,-0.000760838736615588,-0.00484272265898678,-0.00372139381394476,0.0084223245289663,0.00357184743691041,0.00275675734983505,-0.00186573466830275,-0.00211479599145925,0.00761242387006322
"2421",0.00288384687692833,0.0020303457663291,0.00567719679079715,0.0104055619487864,-0.00942272565349944,-0.00293640078489188,-0.00071717938692184,0.00397269608217532,0.00345364201799625,0.0164835036664763
"2422",-0.00515760043778213,0.000506592783606541,-0.00887098386552854,-0.00448899164311867,-0.00266620032521858,-0.00169567274716864,-0.0117224236895006,-0.00256072629578474,0.00492807430938913,0.00810813667656118
"2423",0.0018809335087695,-0.00151889743291322,0.00813683525078801,-0.00636621200819987,0.0059969727241469,0.00160927080295359,0.00290466184154559,-0.000232847136946268,0.000233509767000095,0.0040214617765566
"2424",0.0022439904434397,0.00760676515409209,-0.00484272265898678,0.00934333827268596,0.00158057551590463,0.00178511618769295,-0.00289624921696152,0.00373431988178607,0.00474708949416347,0.0126835420999869
"2425",-0.00146224836903086,-0.00830413183901324,-0.00243306894558803,-0.00555404020045069,-0.00523517618703662,-0.00338575742865277,-0.00726240247133081,-0.00697642582301083,-0.00882968004934037,-0.00329593395865624
"2426",-0.0000456973780924574,0,0.00569097868233404,-0.0132977285756044,0.00843520030274547,0.0022349861538169,0.00512083249820861,-0.00210778755842567,-0.00148473859900955,-0.00925926871340432
"2427",0.00201349051401634,0.00456729280295476,0.000808522205114404,-0.00404308823159705,0.00107149213937885,-0.0000893037035900601,0.00218351687789653,0.00657111833655666,-0.000156495540432733,0.00400528569093561
"2428",-0.00511474545450807,-0.00303097200975255,-0.000807869025068797,0.0027062069080499,-0.00235586425705137,-0.000356584652292491,-0.00484145853711282,-0.00373056546436568,-0.0111146366450433,-0.0119681274213354
"2429",-0.000688713666437302,-0.00430711468522693,-0.00485031695385063,0.000809843647337827,-0.00379444343219182,-0.00160625437017137,0.00364843565428785,0.000468081833877809,-0.000870611077112948,0.00403776877017403
"2430",-0.00188325433964187,-0.00534354409997706,-0.00731113005757034,-0.0086302502180553,-0.00581979964098944,-0.00384356893259385,-0.00933093036042698,-0.0112279585668875,-0.00142596843636289,-0.00335122964418233
"2431",0.00492412765832939,0.0046046820101846,0.00327333007381103,0.00761700081702932,0.0133711206343841,0.00412766499305439,0.0094188166829734,0.00070982408848419,0.00198333989726285,-0.00403491472006745
"2432",-0.00164852722466602,-0.0015278773751648,0,-0.00269963206214296,-0.00385160287577735,-0.0000895305605623786,-0.0016962365606682,-0.00520099759968407,-0.0100554550263946,-0.00945308182100768
"2433",-0.0028439683787973,-0.00178515773026822,0.00163133600801246,-0.0110990785711613,0.00143141297272686,-0.00116186757035874,0.00194221699227004,-0.00166353142207054,-0.00199952013116467,-0.0190865205881448
"2434",0.0000460105482600337,0.00562087054085847,0.0073288394992892,0.00766495756642405,0.00110331596240498,0.00156791534354217,-0.00169636565773923,0.00928348100869036,0.00408720952145547,-0.0111189659261556
"2435",0.0045079102664467,0.0149899206838155,0.00727566875950036,0.0162998820965412,-0.00815651812182883,-0.00259386884650115,0.00800973179531694,0.00117925169915845,0.0102162901251792,0.0112439874393682
"2436",0.00302245124648248,0.0055066019856127,0.00561796470864251,0.0213846385064682,0.00728622555386949,0.00466330934827641,0.00710326796751737,0.0148410157075434,0.0169076953464486,0.00694917489634173
"2437",-0.000091337715093065,-0.000248959210288557,0.00478861486759019,-0.00314060607949462,-0.000716347009670715,0.000535720057762701,0.00573842282326065,-0.00580295030386524,-0.00341856092044179,0.00897172432975935
"2438",-0.0022829535623986,0,-0.00476579331884763,-0.00262512764873257,-0.0125414047877732,-0.0049072305650848,-0.0114110496050166,-0.00256870758656569,-0.00530137973645028,0.0177838964431223
"2439",-0.0239348392693182,-0.0209161378150358,-0.0159616254252044,-0.0336934662592854,-0.0164741215129011,-0.00475198887417361,-0.039797957696538,-0.0255147825606946,-0.00658355691146817,-0.0154570542315235
"2440",0.0143473476178548,0.00890115298939409,0.00811035193900511,0.00681038613873675,0.000516387838425336,0.000900997137109227,0.012146238345554,0.00480425372193283,-0.001262358974359,0
"2441",-0.0143756610361736,-0.019914088996399,-0.0176991460696774,-0.0251624115476015,-0.0113577857167236,-0.00369081220259737,-0.0243722698019667,-0.0207985146194173,-0.00663556384028952,-0.0129693172763443
"2442",-0.000375197831216645,-0.000514495334514309,-0.0065520439634662,0.00305311929690544,0.00149212956517464,0.00225872921477133,0.00304337286974277,-0.00170895611026989,0.00341948310139162,-0.00760708883651384
"2443",0.00999315062246486,0.00797728238558837,0.00494652442731858,0.0171553061071559,-0.00432078884239395,0.000270283686430339,0.00455144696498944,0.00611399733186313,-0.00641937708036144,0.00487798195622902
"2444",-0.00386568750396366,-0.0178708184435823,-0.00820358433658464,-0.00680067968146369,0.00807981539142055,0.00108172343869994,-0.00100691723513002,-0.0110593474261649,-0.00247272068741999,0.00138694364428016
"2445",0.000187336650752545,0.00779833701170252,0.00330854954204374,0.00794292848013511,-0.00326509123343144,-0.00171024556991473,0.00944798720460693,0.00793489386991642,0.002079018104574,-0.00069244007257252
"2446",0.0000470173441911026,0.00206333820365767,0.0140148787192746,0.000543494790867349,0.0034992779977403,0.00153280200355521,-0.00162199575148425,0.00442778115296139,0.000957564634535668,0.00346495601403118
"2447",0.0112454539241151,0.0128701099524231,0.0292683193444581,0.0279741737341372,0.00808732106613674,0.00162046133092386,0.011499598236862,0.00857211213528597,0.0145886078668909,0.0124309117376125
"2448",0.00630145677084881,0.0116901260993136,0.0126381345563149,0.00713313508244195,0.00794873504866422,0.00296645780690152,0.0194023227572044,0.0114133556777394,0.00235721699592717,0.00545709200812983
"2449",-0.00547929428082239,-0.00753595493055881,-0.0140404821098483,-0.0128540097729919,-0.000949114274031659,0.000447863224858347,0.00254571615167132,-0.00408144527788612,0.000627122364192267,-0.0115332945108013
"2450",-0.00810212189224324,-0.0111363548469304,-0.0087026311513686,-0.0146159364462848,0.00635874755153454,0.0028667099799895,0.00117055328905735,0,-0.000783384241545115,0.00686346568920571
"2451",0.00620803345474608,0.000767736603415781,0.0111732650376719,0.0142933693063589,0.00733511600412617,0.00169718447833422,-0.00779537540340924,0.00771447407612724,-0.0072912581585749,-0.00954336553088786
"2452",0.00496348444299533,0.0112533555499574,-0.00157854623374787,0.00904016321940171,-0.00216277180315305,-0.000445923702765749,0.00552421255335256,0.00334933022817396,-0.00315907432098228,0.0233998982825621
"2453",-0.00904712310608102,-0.0144160519769228,-0.00711470992276098,-0.017391345103953,0.00252862913802776,0.000624657939502837,-0.010743587189161,-0.0164522289939346,-0.00118840911750584,0.00605251050862865
"2454",0.00754593641498302,0.0105210771718134,-0.00159220199293086,0.00429076648435722,-0.0089367614632665,-0.00249661225969966,-0.00481297367118139,0.0111515703652236,-0.00341081145395405,0.00334226902923129
"2455",-0.00240419902037381,-0.0015235257188092,-0.00318982132203227,0.00694251052310624,-0.00330031150400256,-0.00232692832720705,-0.0181051643832972,-0.00455530403482884,-0.00254695162804008,0.0086608425336514
"2456",-0.00509747804628857,0.00152585039112307,-0.00559998670126716,-0.0111376219313902,-0.0116954630597766,-0.00457550515011851,-0.0143974643026727,-0.0139692590930305,-0.0347111315033514,-0.0026419718257199
"2457",0.00442510181287625,0.00253925608903294,0.00643607838030191,0.0144810678501628,-0.00465936681570889,-0.00225286094459709,-0.0193491558239017,-0.0134340654728494,-0.0015706538681437,0.00596018324407677
"2458",0.000695416360598333,-0.00607894622013694,-0.00479626978176939,0.000793117151379086,-0.0055725484164787,-0.00207707089818854,0.00169869408796419,-0.0118842318551126,-0.00927301713258011,0.0019750244006882
"2459",-0.0034292167452119,-0.00764519932650454,0,-0.00449040595762129,0.000672475566745545,0.00144789087125985,-0.00143496914151819,-0.00876968281953339,0.000668510758197849,-0.00262808499404299
"2460",0.00520841514603565,0.00231137933535108,0.00321294457740495,0.0108783322451635,-0.00589863006018765,-0.00262109698223656,0.00587852700281499,0,0.00350764996672215,0.011198928205062
"2461",-0.0126297359905929,-0.0148605701018741,-0.00880706088130723,-0.0230972152953798,-0.00225389462550551,-0.000271957408808254,-0.0100001361529047,-0.0171889314508663,-0.00507657273380246,-0.00586324608441957
"2462",0.00131198652739473,-0.00286076982234174,-0.00161552341398208,-0.00188057710350076,0.000978797710992962,0,0.0135119080523329,-0.00154345580457182,0.00158925131938314,-0.00720842462624149
"2463",-0.0032754682313183,-0.00443403052218161,-0.0016181160547396,-0.0088830156201829,0.00376031432954171,0.00208478315212779,0.00556568599139506,0.0108194849563596,0.00242192253920037,0.00660070625287879
"2464",0.000516542946895626,0.00104795810427083,0,0.00162962815027989,-0.0140114751820759,-0.00307532106947739,-0.00334677794708693,-0.00280349806729541,-0.00558192123287449,0.000655728765314612
"2465",-0.00347239848887548,-0.00366421516198645,0.000810401598727362,-0.00108457276699547,0.0063835776622394,0.002177683179859,0.00129158876099877,-0.00536681945906881,0.00268095674697588,0.00131066557908799
"2466",0.00626240335754025,0.0123461006777812,0.00566785189063124,0.0176437963425582,0.00324655859356748,0.0019917068124593,0.00683587474629932,0.0125898648860383,0.00618313836898388,0.00196339129656375
"2467",0.0026672507494887,0.00155661728325573,0.00322064133799782,0.00613488076135904,0.000828227304453533,0.000451599613674469,0.00422783085420719,0.00558248947657924,0.00572997019980015,0.00653165629159558
"2468",-0.0018668599300522,0.00025917074424564,0.00882833079239864,-0.00291606920989806,0.00105287969206969,-0.000903091863339478,-0.00382716851521481,0.00252332671480482,-0.00305509864540421,-0.00908501892228064
"2469",0.000467607933100966,-0.00259012418709259,0,-0.000265995717653622,0.00150278454221531,0.0010849516302216,-0.00128078866976788,-0.00226528440221807,0.000745436487418205,0.00392921932243606
"2470",0.00425262071561683,-0.00129836804460626,0.00159110425844444,0.00425527545179527,-0.00435098629292341,-0.00135477542985907,0.00269292947329669,0.00227042756637053,-0.00223457746859923,0.000652373967855002
"2471",-0.00335041094859378,-0.00260002618303401,0.000794246122462594,0.00105952662299025,0.00263697911850547,-0.000180791894687782,-0.0019182410578279,0.00125832789643976,0.0075481338345742,-0.00456323801298775
"2472",-0.00200776027938832,-0.00547437144167284,-0.00158737921437313,-0.0105820149845479,-0.00676303048235494,-0.00217037040479251,-0.0116590846390477,-0.0103062729953215,-0.00559809001730394,-0.00654883367309145
"2473",-0.00266664584910203,0.00183475815514944,0.0015899029933375,-0.00855614753053668,-0.0108939548545162,-0.00344424839539659,-0.0229454420331365,-0.0111761569295213,0.00182135109014525,0.0059327489710721
"2474",-0.00295565987189239,-0.00130821954003113,0.00158740030322813,-0.00404550291354611,-0.00221826188591334,0.00018168811507735,0.00199004179742612,-0.00616475208154399,0.00471035443830492,-0.00655305811402018
"2475",0.0000471342157475352,-0.00104784282369175,0.0007923580068534,0.0056864747327996,0.00613286665331803,0.000818837990992582,0.0148307896004547,0.00749527514614567,0.00296101327585108,-0.0131925678921104
"2476",-0.00724536253600916,-0.00445856586976356,-0.00395896894499981,-0.00807743955302287,0.0000760304627447361,0.0000361395076220461,-0.0220513708319905,-0.00384807277934451,0.00647860412533041,0.00467914912177814
"2477",-0.00601860252229691,-0.00711277778487773,-0.00635918952566294,-0.0119434304052429,0.00435121104745018,0.00300213139370609,-0.0128084265246907,0.000772378132541052,0.00741461727170334,-0.011976089318696
"2478",-0.00457724324954434,-0.0021224920765549,0.00239989408630681,-0.00274745485220673,-0.00767623266949324,-0.000634810732857649,-0.00581153998172868,0.00257345676614862,0.0053381106869792,-0.00336702670285538
"2479",-0.00110137929486009,-0.0090403046697155,-0.0119711448455531,-0.0101928334653643,0.00896059792067283,0.00308614174701938,0.00530172963015918,-0.00770025977644295,0.000724022508671984,-0.00675673420271494
"2480",0.02205675194794,0.0160987306482849,0.007067796886286,0.0361814463486601,-0.008501919794068,-0.00416248676141207,0.0163625754717327,0.00931202325161595,-0.0180078544738954,0.00408164694177549
"2481",0.00450394144179223,0.00316886716477427,-0.00120309639231997,0.00644643535599121,-0.00405703187388529,-0.00354368687375517,0.00612026786939079,0.00256267615162997,-0.0041752189246792,-0.00135499503103398
"2482",0.010602203474694,0.00500134286684317,-0.00843211777843456,-0.0325594726249419,-0.0424322319805887,-0.0152289498142567,-0.0185135457823911,-0.00434550125429056,-0.000657686621651554,0.00474898719275374
"2483",0.00249544997536755,-0.00366674856166804,0.000809995506815708,-0.0284137164936527,-0.0147707204585984,-0.00601929162596859,-0.0181894428229691,-0.0269579099066729,-0.0148897501627139,-0.00810266141648341
"2484",-0.00230488840821275,-0.00972678224885215,0.00141610299859818,-0.0190233215188182,-0.00562222607095253,-0.00204921094077148,0.00535205642999892,-0.00765131197336766,-0.0221294530271399,-0.0190606052729353
"2485",0.000785451305220786,-0.0082292863702822,0.00121219656033267,-0.0072358120129743,-0.00598169452868991,-0.00578802213782392,0.0169261114782746,-0.0124965570244908,-0.0084542870786386,-0.00208185917709702
"2486",0.00780276818525283,0.00588867460786324,0.0016142194400377,0.0201166437499278,0.00494579625837321,0,-0.00362428648420865,0.00700028518350093,0.00869866498407834,0.0222531114282418
"2487",-0.00187824028611006,-0.0119745195932006,-0.00483485380511139,-0.00828807021708278,0.00902330097789172,0.00093903095999992,-0.00215540287511362,-0.0131016730701958,-0.00298843913110214,-0.0122448708106266
"2488",0.00514068218958919,0.00457852786953694,0.0149798054214234,0.00144098150397109,-0.0147143213135938,-0.00440915732321745,-0.00823563918812775,0.0149009245627292,-0.00513829763993223,0.00206601655464245
"2489",-0.00223758017901077,-0.0109920081903816,-0.0149582825618577,-0.0046045807107481,-0.00288782418421973,-0.00442853269113563,0.00299495667940675,-0.0085419448102152,-0.00878020158010162,0.0082475228783081
"2490",0.00755140162802381,0.00975890952754099,0.00809885754243034,0.00982963644135126,0.00248279268792229,0.000852060643773411,0.000135820290106947,0.00215356815117729,0.00373425959645224,0.0279482321863713
"2491",0.00195329114274934,0.0010737223278694,0.0024100802617204,0.0151731823314931,-0.00033043767308083,0.000945609547320814,0.0170984685478077,0.00537352825905768,-0.000346089282815432,-0.00132631000327676
"2492",0.000544013604544702,-0.0072404863779717,0,-0.0107161969996484,-0.00388064052743209,-0.00359009972462132,-0.0054700806827932,-0.00213772619742114,-0.0198199842494375,0.00398407763104802
"2493",0.00371544065277551,0.00810378146257595,-0.00841513851374687,0.0048458880349993,0.00149210603860928,-0.000853128287876315,0.00509777259544664,0.00133903898129062,-0.00565120529801322,-0.00727510080633487
"2494",-0.00469494549352489,-0.0112542053455486,0.00868852025258904,0.00397172123160461,0.00736613184142909,0.00455465480559347,0.00347051812540955,0.00748860437156118,0.0105674628312986,0.00333106690960094
"2495",0.00195022681532775,0.00840124719349267,0.00100168627622743,0.00141267212497809,0.00419036476488444,0.00103951184208206,0.00824657980676746,0.0039818922667576,-0.00465734609866397,-0.0199203198141998
"2496",-0.00239893515800838,-0.00080611308483225,-0.00160095386365633,0.00169311506731318,-0.0162004163256466,-0.00670063326786585,-0.0125326708660924,0.000264435758688286,-0.0134192375762137,0.0304878065787826
"2497",-0.00367560156377389,-0.00134504952539805,-0.00841844810814474,-0.0118308563777816,-0.0105585065096747,-0.0038146510291962,-0.0157647523027716,-0.0129526169549385,-0.00187918568232659,0.0184088928598929
"2498",0.00050096411460121,0.0029627981907856,0.00303211430700312,0.00114013074727692,0.00732744251551165,0.0044883843164909,0.0105873783525647,0.0072309329844944,0.00537921816945297,0.00710139187360448
"2499",0.00600885181234934,0.0158430586950693,-0.00120909367134381,0.00825742224405102,-0.00108682008507788,-0.000380190686212978,0.00792515484423451,0.00451989973974243,-0.00535043700151983,0.00512820106818124
"2500",0.00316742213891863,0.00978054477025436,0.00443891044348366,0.00536589399916698,-0.000753259097910131,0.000380335286146449,0.0063961822762939,0.00608799107929503,-0.00098620225043744,-0.00446429040277008
"2501",0.0130807265578898,0.0141361795103181,0.0148655216547371,0.016853740206477,0.00854415699506617,0.00332783804023218,0.0194652535992548,0.0142068469643066,0.0035897155164677,-0.0076874068323729
"2502",0.00244872398394369,-0.0043882478091134,0.0114805365683655,0.00441984388323546,-0.0117942433956341,-0.00379022922183891,0.00506541316631615,-0.000778317678383544,-0.00232497536752252,0.00193683988393856
"2503",0.00604047354444859,0.00518530702376729,0.00293545770326764,-0.00522557698395609,-0.0124390540319584,-0.00513665154643694,-0.00077535437319487,0.000778923928647313,-0.0104866720444563,0.0051545684159735
"2504",-0.0011478412233179,-0.0015476100557229,-0.00975616473538754,-0.00663526532740355,0.00187234493792499,0.000191249461676257,0.00620813236064244,-0.00544756463221918,0.00380432964122579,0.00641030081676885
"2505",0.00667409219156978,0.011624881770014,0.0118225998887822,0.0111328850754264,0.0035677579849791,0.000573393270020039,0,0.00808569666097081,-0.00333877458942422,0.00254773579355727
"2506",-0.00825434015552451,-0.0145556632179705,-0.0153844972427879,-0.0297276510480933,-0.0111732850903969,-0.00831162479727587,-0.0185090502228461,-0.0165589690347874,-0.0146672253870682,-0.00952992615734338
"2507",0.00411721042537661,-0.000259009857141002,0,0.00170233326853575,0.00505084188938887,-0.00279405771543806,-0.00746469536976113,-0.0144701948306275,-0.013691132708056,-0.00128285619031576
"2508",-0.00195588431774019,0.0031103207068246,-0.0087026311513686,-0.00453133898924696,-0.00229962915844317,0.0012559474619287,0.0133266317780192,0.000739579498844067,0.00661456145386863,0.00449589628991709
"2509",0.00217737429817388,-0.0036174797307349,0.00857937101521333,-0.00682793280413396,0.0107564155674695,0.00463134888703332,0.0110677389768699,0,0.00499762133278225,-0.00575452855061109
"2510",0.00385768641258344,0.00363061340112347,0.000989223359052493,0.0034373593216559,-0.00498330093412247,-0.00211265523459192,0.00180273229778249,0.00653393625840182,-0.00736711510699384,0.00450167871434171
"2511",-0.00278270933099201,0.00155038094225879,-0.00533814874620586,-0.00415763230108601,0.00441405123638572,0.00163627186528958,-0.0123055245406665,0.000282253221779216,0.000556610069982311,-0.00576196249489347
"2512",-0.00172757576983273,-0.00179365080311122,-0.0016080689218011,-0.0118875843928827,-0.00178794565574492,-0.000433334975470046,-0.00184770619625585,-0.00395019446179068,-0.00241077426816461,-0.00128774623731354
"2513",0.00146436676670736,0.00286456900604581,0.00181188029469825,0.00586845449117535,0.00203702173085452,0.000962829951520972,0.00264429316960912,0.00481577209037964,0.00316018229055426,0.00193420953618118
"2514",0.00248113185746091,0.00129848645526942,-0.00622978850052258,0.00437589709957065,-0.00321893800776563,-0.00144297384104475,0.00118699584696058,0.00535656138832374,0.00583709811915112,0.015444003425422
"2515",-0.00826460261205209,-0.00622414269811666,-0.00141551688143693,0.00755131276155319,0.00730871189490645,0.00366089712297835,-0.00592707324574493,-0.0070106180074756,0.00276347646948194,0.000633704922959666
"2516",-0.000222837377038987,0.00704599457521748,-0.0101255988208752,0.0164313849511095,0.00354332355307574,0.00307111198579713,0.00993742402727515,0.0104489306455475,0.0131361380384334,0.00126673755373652
"2517",-0.00365494224781038,0.00570092973534786,-0.000409140361173121,-0.00709021535865395,0.00151332250917346,0.00296588702122236,0.00944630597306118,0.0083847672294397,-0.00616556345846808,0.0018974420434541
"2518",0.00765008915940579,0.00231906770749335,0.0081866295744395,0.0119965726440947,0.00428113181937295,-0.00047665453904211,0.00402909274495888,0.000831240244102416,0.00784599938102359,-0.0119949157764663
"2519",0.00594916012144897,0.00874022816271225,0.0200973794707395,0.00762080112462349,0.00384488464766775,0.00114516677704857,0.0137219377888027,0.010523744918618,0.00353037020430547,0.00766769250680732
"2520",-0.000794446301255469,0.0086647767071828,0.00577122146174802,0.0109242761796342,0.0156533906383589,0.00648318602284559,0.00344779937331996,0.0150725435546564,0.0155150729251752,0.00507298460463712
"2521",0.00357771673789964,-0.00429517165032223,-0.00158307836347038,-0.00415628647354194,-0.00918176068048515,-0.00454702752888014,-0.00216349851921238,-0.000270210062075282,-0.00737255272033122,-0.00126187729913718
"2522",-0.00330068745062539,-0.00380622194144142,0.000991083888692623,-0.000834726657825358,0.00802566535617744,0.00380641655835379,-0.00663181409954983,-0.00189024206186761,0.00823264429530202,-0.0151611396094232
"2523",0,0,-0.00376170351730831,0.00584784861520915,-0.000656581554552393,-0.000473778906949662,-0.00937209726569777,-0.000541363995198552,0.00426026456483997,-0.00448993064839287
"2524",0.00282587402697509,0.00534901484814365,0.00655814060505455,0.0119048329426903,0.00336770273186926,0.00113819379109326,-0.00427684234086978,-0.00243602047375835,0.00309322133286405,0.0109535241994081
"2525",-0.00250987461292684,0.00177349993215992,-0.00157941201118128,0.00437761535614389,-0.00221038832249476,0.00056826272126731,0.00455543285809012,-0.00407055288326141,0.0036123700440529,0.0146590152638848
"2526",0.00229537265313184,0.00379359743935348,0.00632768355008784,-0.000817218078311588,-0.00475844144564685,-0.00217763243083713,-0.00103637958066471,-0.00108997584325143,0.00263361416438879,-0.00188439640516536
"2527",-0.00352340036613308,-0.000755846587652598,-0.0112006175049303,-0.000545335604600461,0.0104692017611592,0.00502879890115371,0.00674447918542409,0.000272718081644863,0.0143595045474083,-0.000629382790976241
"2528",0.00221003516103413,-0.00378211914845306,-0.000198642955844042,-0.00545551257239241,-0.0128079372329855,-0.00708078698175663,0.00167466541288386,0.000545352515879172,-0.00845917148828956,-0.008816065726727
"2529",-0.00370452229974694,-0.00253099446464655,-0.00278286955724194,-0.00301697350156638,-0.00685901165485747,-0.0038032868016441,-0.010418085846074,-0.00981180767105139,-0.000870601526840709,-0.00317664205244783
"2530",0.00367392920517062,0.00532846138402343,0.00637842796997545,0.0019256483845167,-0.00199692305585197,0.000476881846938948,0.00636863162832202,0.00385348919611417,0.00243971427480294,0.0114722499988849
"2531",-0.00260227483046038,0.00328137031188236,0.000594088797734704,0.0148270569749624,0.0100049909433235,0.00524744858693982,0.00761989883101477,0.00795159795073253,0.00643196854153927,0
"2532",0.00641192069678653,0.00201254826811592,0.00257336232983607,0.0062229211077367,-0.0068518476802224,-0.00379607770766222,0.00230703850678848,0.00108819705190211,-0.00449092318429123,0.00252050941723025
"2533",0.00865551118260455,0.0120511733746524,0.0104639001615463,0.0110244592132693,-0.0125505010042011,-0.00495390406586704,-0.00537098560592064,0.000543426042516337,-0.00824149409841668,-0.00628526933019513
"2534",-0.00104530482878629,-0.00620192319802526,0.00136766917038544,-0.00425536829860129,0.00336683800293636,0.00134033752256624,-0.00102826995030203,-0.00461700135763288,-0.009272200839748,0.00442745156679414
"2535",-0.00156983936953636,-0.000499243626010948,-0.00819507373889461,0.000801398748848881,0.0036073408826891,0.00124311114177589,-0.009395128921871,-0.00136412539642139,0.00203069041090065,-0.00818635137568224
"2536",-0.00620176026995189,-0.00874131828248248,-0.00275431775039814,-0.00533757885371866,-0.0030093504941775,-0.00028656348497913,-0.00688565718933232,-0.00109295398804843,0.00422947403699836,-0.00571427301828686
"2537",-0.0000877447645776241,0.00377917792158833,-0.00236716587615005,0.00187834439384749,0.00695927678084818,0.00343866619063449,0.007849036402507,0.00957323196488957,0.0138633147857918,0.00574711359443247
"2538",0.000395421879109126,0.00326325038439301,0.00533898429387358,0.000535351875829315,-0.00618336796058461,-0.00191634048718048,-0.0118118875594656,0.00189638742332776,-0.00302904362538192,0.0107936340731034
"2539",0.000658919415098991,-0.00100095402576972,-0.000393367056473082,0.00428281959216603,-0.000419821657313912,0.000382101265646195,0.0111651186845563,-0.00243374021693377,0.00555554701967576,0
"2540",0.00689306532363032,0.0040070894933697,0.00452573907890552,0.00612992666580281,-0.000419780144993664,0.000763778274778915,0.00675489105645277,0.00542168218861572,0.00250346175771621,-0.000628132135055082
"2541",-0.001787817673089,-0.00947872216163737,-0.0015670985090328,-0.00238411216811607,0.00605020935167411,0.00477045683397326,-0.00335483485716837,-0.00188740918955965,0.0135193321325926,-0.00628526933019513
"2542",0.0000437172102030203,-0.00125902747056506,-0.000588638418962173,-0.00504507797170339,0.0073505528095883,0.00180442996670105,-0.00142406518786775,0.00216091543931229,-0.00203906547253352,-0.00442764686394759
"2543",0.0013103846925393,0.00252153205859806,0.00294467809241827,0.00613822140535336,0.013598803707106,0.00407568998480334,0.00726040357045532,0.00539089711437257,0.00621490725536278,0.00381195738522355
"2544",0.00593259105414901,0.00402391944384473,-0.00137007854487714,0.0045093712544626,-0.0115347474536788,-0.00594686571239511,0.00308918934808156,0.00428942023602374,-0.00761486576504167,0.0050632218761828
"2545",0.00394618218828069,0,0.00705605879750415,0.00924212936540303,-0.000579395860808574,-0.000665069146421171,0.00769928244374385,0.00106792618797336,0.00264299597030426,0.0107053384040592
"2546",0.0054427099283505,0.0045089784226362,0.0038926346481678,0.00313972526534179,-0.00314701042197341,-0.00152066305376009,0.00331084687230998,-0.00293321077133191,-0.00680267868712037,-0.0112149924655612
"2547",0.00399531217314886,0.000748336411536821,-0.00717354722988917,0.00104333670624057,-0.00722690948271076,-0.00361655496898972,-0.00558439924195642,0.000267457385086045,0.00111298798511172,0.00126028713508397
"2548",0.00522027846356843,0.00274107749348462,-0.000976179084352213,0.00807695702322619,-0.00460184265387809,-0.00191039428403483,-0.000893659771184829,0.00187173299152521,0.00444707944924305,0.00125863603933829
"2549",-0.000851234367105991,0.00472165339998631,0.0011726581030711,-0.00361836771855262,0.00546366699282075,0.00401970686387476,0.00472666689117363,0.000800436136135341,0.00536402738264852,-0.00628526933019513
"2550",0.00157628852865543,-0.00321562893528105,-0.00058560126906182,-0.00415050131909678,0.00593596241106709,0.00266891643068323,0.0016530614692436,-0.00106678693826512,-0.0033875507556308,-0.00189763734060744
"2551",0.00595517372264642,0.00124089317216436,0.00840010990280105,0.0109404604500907,-0.00174521431805508,-0.000475343533529071,0.0125665565644317,-0.00240255527811739,0.000594833446634802,-0.00126734462309919
"2552",-0.000888037909210548,0,0.00116237104316563,0.0030918835432161,0.00166493157201053,0.00161660192047153,-0.00250737897997322,0.00240834145158342,0.00135884501061567,-0.00507620312805912
"2553",0.000677126376396719,0.00272602417953638,-0.000967606015941369,0.000256826045995195,0.00299227454620365,0.0026590229852177,0.00427314785577559,0.00453840765406444,0.00873545895223615,0.00318873197427805
"2554",0.00126895379814229,-0.00889773331518162,-0.00213046534719108,-0.0118130025310037,0.0111047964752546,0.00464059889104518,0.00500574817128863,-0.00212607599588366,0.00638973421238043,-0.00190709233946518
"2555",0.00156284324533473,0.00174563728176347,-0.00310560456499609,-0.00311862243565053,-0.00590108417176605,-0.0035822715931052,0.0052295511163678,-0.0039945444088324,-0.00484539694683539,-0.00254780134871879
"2556",-0.00269922187852611,-0.00174259534236676,-0.00253119263241841,-0.00964530310053924,0.00370991402959242,-0.000473050087338223,-0.00396377869017817,0,0.000923438526105436,0.00383143097049166
"2557",0.013997544476545,0.0117208513778566,0.011711932645359,0.0155304035325612,-0.0167561404143637,-0.0069664737322449,-0.00310900993659491,0.000802189508483986,-0.00142585755030133,0.00445286527660071
"2558",-0.00629738726995732,-0.0036973925215037,-0.00945396507770557,-0.0176257193461409,-0.003599336798363,-0.0028636102091244,-0.00411676677005723,-0.0125568078166178,-0.0124306738187582,-0.0158327854283856
"2559",0.000629601603776786,0.00841174127417554,0.000584232424516884,0.00765158312162728,0.002604205288947,0.000957566817019861,-0.00237995119025658,0.00405850320230372,-0.000595339333299139,0.0051480673719293
"2560",-0.00297793578731897,-0.00515197933218881,-0.00233597423016452,0.000523773546083239,-0.00477565165141025,-0.000191521602316946,-0.00464615974657034,-0.00161675575512177,-0.00672284049488825,-0.00128045807361343
"2561",-0.0029869737039705,-0.00567208589159396,-0.00234144378250178,0.00104677419273358,-0.00303107447186834,-0.00143489962257004,-0.00428910768580171,-0.00485854022918186,-0.00805347834087144,-0.00448725015697193
"2562",-0.00185657199752809,-0.00421626074793802,-0.00312929310750232,-0.00941167710692248,-0.00540466520569627,-0.00335204319919824,-0.0153300232978704,-0.00867911835488477,-0.00621869931092334,-0.0225369177448197
"2563",0.00126824262216241,0.00797007402280592,0,-0.00791767631638118,-0.00798073117033782,-0.00278699648902048,-0.0127379498105936,0.000547371528188068,-0.0051277334456411,-0.00856391818071489
"2564",0.00350408421226756,0.00889542587552472,0.00725925545124384,0.011173212724702,0.00350915915433747,0.002120063583126,-0.00247622126604929,0.000273454487948355,0.00218397831585593,-0.00930240351013967
"2565",0.000504967747655627,0.0039187624701662,0.00506413214011769,0.0139437810553684,-0.00631144812149054,-0.00250046738784948,0.00156791149128366,0.00191346245000745,0.000174311365286783,-0.00134129435353814
"2566",-0.00382667477613463,-0.00731890831984305,-0.00697660464156658,-0.00570837810110747,0.00480653038543233,0.00106051781121441,-0.000913346232412349,-0.00818546845485246,-0.00540347752141324,-0.00402956400638621
"2567",0.00865346427644575,0.0135169545735745,0.0101482766939005,0.0260959108673648,0.0122149102925839,0.00876446895663108,0.0184098760670601,0.0159560901169946,0.0186645368384717,0.00876603378785168
"2568",-0.00196679238728203,0.0104267189554459,-0.00193213992819286,0.00610375241894068,-0.00506341894665796,-0.00276902272115742,-0.00166672196681106,0.0119140610741635,0.00412905806451613,-0.00133694889041081
"2569",-0.00175628623922197,0.00191963418032004,0.00329092332896663,-0.00176939639504703,0.00627665346892248,0.00268080497575318,0.00423773217401036,0.00263648667465266,0.0022273193979101,0.00334674345417874
"2570",-0.00109680203397067,-0.00191595624522367,0.000192916551013722,0.0116485841285048,0.0042987058848587,0.00238707354792367,-0.00038382170549589,0.000804988867886491,0.00444485861090449,-0.000667102292611355
"2571",-0.0128396254567116,-0.00359978898565694,-0.00771610592965055,-0.0110138657863131,0.00830883642509939,0.00333398922866879,-0.0031978719996949,-0.0075067408605104,0.00876520281226778,-0.00534051833327187
"2572",0.00235316658674178,0,0.00136083816258492,0.00480895759237554,0.00399545941916934,0.00189871800113472,0.000513261357844241,0.0027014167757855,0.00244643999960825,-0.000671062731966487
"2573",-0.00106693896534815,0.00120424723030488,0.000776582510718882,0.000251817771555141,-0.0014098156166964,-0.00104217708703658,0.00743967023452163,0.00404076064475722,-0.00134649497018424,-0.00201488568513231
"2574",-0.000726570081885924,0.00360844881822842,0.00620753347389047,0.00251840786784929,0.003570196530573,0.000569225007692742,-0.000707035457979899,0.00295172136254651,0.00160110392855994,0.00336476113458128
"2575",-0.00102624490080683,0.00527311868793201,0.000578424903030283,-0.00276320337007108,0.00454992670454235,0.00246491872838206,-0.00681728599172537,-0.000535238559549511,0.00563686685481346,-0.00134129435353814
"2576",0.00727683322865791,0.00023843231029308,0.00847779050997111,0.00277085981926151,-0.00667028943947512,-0.00340469169968505,0.00440338505552007,-0.000802700208162754,-0.00409937257675375,0.00604431144893303
"2577",0.000934848081634465,-0.000953423816419052,-0.00133735785228317,0.00175828460679561,0.00596907511322753,0.00284680128581272,0.00438418030198373,0.00267856912971243,0.00243616429405091,0.00934580402420737
"2578",0.00318424345690382,-0.00381788187884613,-0.00554824950578392,-0.00526581051277752,-0.0080764818165302,-0.00283872001402663,0.00295291036624268,-0.00534358797024104,-0.0072069134801489,0.00396826774429404
"2579",-0.00232760000833565,0.00239530488338602,-0.009234243994378,-0.00705828412172327,0.00290788998354463,0.00199272553168406,0.00473623764313547,0.0045665689340979,0.00211023886122863,0.00197625751826047
"2580",-0.00173928836426529,-0.00382314715306309,0.00504856245789309,0.005585115599686,0.0100868951300916,0.00492269566694903,0.000891991671073233,-0.00106965091891176,0.0053065784593449,-0.00394485458956617
"2581",0.00063725119751723,0.00143906781298697,-0.00347751898115156,0.0005051047989586,-0.00542457751624892,-0.00141586408660166,-0.000891196731011901,0.00214137026607597,0.0022622958066576,0.00990112731437764
"2582",-0.00297238472389372,-0.00670635680364251,-0.00697961417527004,-0.00302812469026936,0.003057280604287,0.00189042176690291,0.000254885020888329,-0.00160241371171721,0,0.00196069013709699
"2583",0.00281120669829771,0.00337593631499433,-0.00507607934606946,-0.00177174407320924,-0.00148278328093321,-0.000660382132687931,0.00687815146792459,0.00909575411798946,-0.00367833965026731,0.00260929445926572
"2584",-0.00101963685707351,-0.00144214929942332,0.00215862008465884,-0.00177477996801234,-0.00404273002357236,-0.00302097072468743,0.00113865379477773,0,0.00234937909045141,0.00260250376062299
"2585",0.00059538022964345,-0.000962602424151027,-0.00234977849809492,-0.00406405470104532,0.0046390834084431,0.00179912266291171,0.00694946284429721,-0.00397695711016866,0,0.00778704458108392
"2586",-0.00118977264711828,0.00602260777388453,0.005102916886631,-0.00229531137595762,0.00948286736333603,0.00463156448385704,0.00552148739241543,0.00904988394114525,0.0144818601580603,0.00193185131067319
"2587",-0.00438179560405416,-0.00119730016460229,-0.00331953410031871,0.00485687223381781,0.00547303244111874,0.00310477274528842,-0.00224629573928015,0.00580352936868067,0.00684870852630226,0
"2588",-0.00649501135743358,-0.00695274391045941,-0.00842471471963524,-0.00432457389914864,0.00308714042240155,0.00300097094078722,-0.00200133045897133,-0.0020985000764302,0.00475332744025558,0.00321332361178372
"2589",0.00885985025495395,0.00627714605303065,0.0106696964283806,0.0104750972642398,-0.00307763931765848,-0.00158968252076741,0.0125331106195241,0.0113010564835776,-0.00293637851445971,-0.00576545622459146
"2590",-0.0029842634088022,-0.00527828451928669,-0.00312792601824285,-0.0126423033537344,0.0130798984001015,0.00571337423900875,0.00235186182224667,0.000519814821712927,0.00474478083679286,-0.00386605894290903
"2591",-0.00183854861629096,-0.00337682983485821,-0.000588407500659582,-0.00614568124507953,-0.00545295831716142,-0.00260766002111623,-0.00160561120997105,-0.00831185309442883,-0.00887475166910923,-0.0174644522676406
"2592",0.00813917894131433,0.00774458271198109,0.00608333701858621,0.0123678657302932,-0.00387057090925247,-0.00224090712638458,0.000618509539508816,0.00392898079498871,0.00188939451517145,-0.00394991328905014
"2593",-0.00318695376026734,0.000240254970751641,0.00370579830383289,0,0,0.000468091578306851,-0.00395554843296653,-0.00495705464799445,0.00286978519899783,-0.00991407848530956
"2594",0.0109979221564875,0.0362543990727437,0.0069956452875235,0.0142528805525413,-0.00493751063823911,-0.00205754330369856,-0.00868704717253677,0.00498174945227192,-0.00678599471483921,-0.00333780678179185
"2595",0.00581858699768523,0.00880449334264033,0.0036665275893617,0.00878303061256203,-0.0120395301324693,-0.0051552859984304,0.00287924907763304,0.00417423472053891,-0.0101251479224939,0.00468855149106728
"2596",-0.000628716122163531,-0.00390452220996029,0.00115365505637066,-0.00373135263953883,0.00551681542575233,0.00263773332189032,-0.00661590538861012,-0.00363729567264037,0.00490641164241157,-0.00533332912498308
"2597",0.000838839255357771,0.000691712010259637,0.000768331451396431,-0.0012484068936307,-0.000327637919719015,0.00065785586228384,0.00113095909403405,0.00130398855767377,-0.00372390776974207,-0.00536192604130525
"2598",-0.00217924118577906,-0.00115215708641392,-0.00479764387472803,0.00149989649507831,0.0022116240251322,0.00103305393156194,-0.00928817213470468,-0.00572956474194641,0.00315639175310567,-0.0026954503170562
"2599",0.00251997574656548,0.00392163608598328,0.0038565853640351,0.00574126001337727,-0.00831306099492546,-0.00216061916796262,0.00608136917962465,0,-0.00910821418667418,0.00202706893995463
"2600",0.000377080191859003,0.00689335437167027,0.00307333064143367,0.00719801280754484,0.00512063709670563,0.00207096381796013,-0.00251859434360369,0.0112625768705021,-0.000167092841432237,-0.0107889326307644
"2601",-0.00121448198497376,-0.00251025667206284,0.00248936617333029,-0.00665354066462209,0.000657384601531197,-0.0020666837906067,-0.0119936768840041,-0.00466181295744772,-0.0139573670880507,-0.00408999375384422
"2602",0.00117417398486008,0.0148707412700237,0.00248332510321436,-0.0111635113175481,-0.00492703965550267,-0.00225988118867693,-0.00434440632725241,-0.00208184056640992,-0.0100864720269586,-0.0239561487734999
"2603",0.00393694265534328,0.0114967950229403,0.00552590843140677,0.0082789976501676,0.000907807058279753,0.000188573821060523,0.00962536983042805,0.00573666473366297,0.00188373146773069,0.0140251252850372
"2604",-0.00016681906006466,-0.0104746457932766,0.000379139419816266,-0.000248747597336507,-0.00544157453615668,-0.00245272038823308,-0.0057201209479677,0,-0.00222204935950687,-0.00414932118355293
"2605",-0.000918056010227986,-0.000225221852377167,-0.00322039892211023,0.012692806670304,-0.0000827973569587082,-0.00113521600262945,-0.00536958722032377,-0.00103708056805452,-0.00599569164882219,-0.00486111622344032
"2606",0.00179584551207368,0.00270309889390408,-0.00456096508161852,0.00663544847801134,-0.00116064795489701,-0.00037865444109908,0.00539857534148536,0.00103815722073475,-0.0000861869861390474,0.0160502406843015
"2607",-0.00204267749214504,-0.00292040355568213,-0.00267273324085981,0.00219727141567994,0,0.000758058360095015,-0.00536958722032377,0.000518386460151676,0.00396414164112247,0.0041208935885988
"2608",-0.0016711512276566,0.00788621818787094,0.002488493427939,0.00414137165738016,0.00755296914133963,0.00511090262046832,-0.00269940875751384,0.00181378154803613,0.00283263519313293,0
"2609",0.00552360691444131,0.00581281152505864,0.00286425112387723,0.010189150448878,-0.00271845328115006,-0.000659210893546591,0.00360916797887212,0.00517327150829638,0.00265340233410249,0.00547195189069516
"2610",-0.000915610955030344,0.0102244380615419,0.00076158815866556,0.000960857668476978,0.00371714453975325,0.00131913140421469,-0.00565064947406713,0.000257533857732639,0.00435379037351713,0.00136059565705837
"2611",-0.01774397899923,-0.0138613231578141,-0.00152215709143322,-0.0170346581617168,0.0145668945072592,0.00799937029841358,0.00529519212494645,-0.0036017372007886,0.0181895364523665,0.00679338516144568
"2612",0.00402855097791233,0.00133869235760731,0.00266772066206955,-0.0165977262744018,0.00113539558359244,-0.00028018719402878,0.00269790728370611,-0.00335651155889383,-0.00818100836312718,-0.00269901859172683
"2613",0.00650407981935031,0.0131461891803255,0.00817174907096829,0.0213453758787325,0.00234969841702437,-0.000279809633472627,0.00589349983911536,0.00595859445009927,0.00496594571106734,0.0196211203497609
"2614",0.00507744075907657,0.00241916512798546,-0.000565558928756871,0.000971986489439747,-0.00274820864269243,-0.00112129731381749,0.00292968969194463,0.00103001422205584,0.00418760461997314,0.00663567772410345
"2615",0.00221280589363038,-0.00153585800142664,0.00132036443976702,0.000971355048884126,-0.00672789092852821,-0.00261833762100894,0.00228594945006777,-0.00205793929614839,-0.00633864042804599,-0.00329593395865624
"2616",0.0023328564813232,0.00153822048967367,-0.00150690202328696,0.00388060941339075,0.00563079779145981,0.00206248968546108,0.00671577527069922,0.00386685723600899,0.00394495554763252,-0.00198416790706935
"2617",0.00477935397050411,-0.000877588658384054,0.00264104844718038,0.00483195880580767,0.000324550364839471,0.00056156340635205,0.00213962546691926,0.000256882806071834,-0.0010868489165885,-0.0218687617841493
"2618",-0.000206747050329081,-0.00483096524461157,0.000564356441123515,0.00360674870331823,0.001703737361475,0.000654787946722912,-0.0061543078651709,0.00154029171284997,0.00887176074141882,0.00745254240077342
"2619",-0.000868780321898077,-0.00154457291633758,0.00206864685733166,-0.00527077086957162,0.00494009375404603,0.00252305647752982,-0.00391751065819601,0,-0.00331841709541714,-0.00806996786866232
"2620",-0.000248429381559223,0.00309390049654845,0,-0.00770701086025938,0.00249824848338709,0.000466433993695947,0.000253606913642734,0.0030762107393556,0.003995372099179,-0.0108473798076169
"2621",0.00795223375114529,0.00638914542359648,0.00900724155297561,0.00849502730933982,0.000104599034631114,-0.000522674568324888,0.00405880451115248,0.00920014811695657,0.000829033307186977,-0.00685405688185781
"2622",0.00332845338129917,0.00656737479486802,0.021015336472177,0.00505426763831496,0.0118404064744313,0.00438842112146909,0.00985367834526918,0.00734341218952506,0.00737243201315074,-0.0048309230214546
"2623",-0.00073713840340639,-0.00587207795883682,-0.00382510462257657,-0.00119749208412412,-0.00620920713466333,-0.00167354419334498,-0.00312755732845338,-0.00276529748969279,0.000986777395059812,-0.00554777457712019
"2624",-0.00319700945552703,-0.00371909064967268,0.000731350574751932,0.000479571116265065,0.00544712668143066,0.00316616290890193,-0.00501949100584365,-0.00151209703049338,0.0112543741578648,0.00697340510093514
"2625",0.00185041450998003,-0.000219583880515017,-0.0003654080459915,-0.00119804473795015,-0.0047802194888954,-0.00185672106012791,0.00416214298310291,0.00403922391564215,-0.00528026816052429,-0.0138503695092584
"2626",0.000492449817042884,-0.00373376981907603,-0.00237606852510197,0.00599782048993647,-0.00264166950231925,-0.0015806803807763,-0.00163282839474954,-0.00402297422195286,-0.0065332382164125,0
"2627",-0.00151770299082898,-0.00286613471300101,-0.00897776394559013,-0.00763154870963623,-0.00152482266514298,-0.000931490823722236,0.00641603777717714,-0.00732161385020569,-0.00912454567818255,0.00561797306157019
"2628",-0.000205541519569974,-0.00508499660352491,0.00314298083347109,-0.00528723774775308,-0.000321602114201958,-0.000186248501734765,0.00662480692031298,0.000254400241471942,-0.00149328022653661,-0.0090782320655145
"2629",0.00489005371405948,0.00577764262029734,0.00552892691490992,0.00483195880580767,0.000160814008262511,0.000372793748855793,0.00211123385491852,0.00991621982205526,0.000997025581613187,0.00422841721504996
"2630",-0.00126779256362164,-0.00176753891338044,-0.000549829488926901,-0.000240477415349605,0.0154366016955072,0.00522005290664929,0.00322173280630089,0.00251736683178461,-0.00547811241339369,-0.0175439077995795
"2631",-0.00192420520668546,-0.00996020442049483,-0.00971943481584525,-0.0103414687737421,-0.00158348102816375,-0.00176190379388153,0.00345830363858024,-0.00502235940903972,-0.00417292605575026,0.00428580271427803
"2632",0.000218445041467952,0.0111782095723296,0.00407403975198628,0.00170113270823391,0.00198242465609666,0.000557312069756621,-0.000615226616610287,0.00349108798607323,0.000167582970164393,0.00426729339038379
"2633",0.00832509401363501,0.00375872868494964,0.00313538684817538,0.00994651446528771,-0.00142475991782642,-0.00278538222182234,0.00172424647758862,-0.00126976662826495,-0.00762523906905432,-0.00637392368741607
"2634",-0.00674408488087042,-0.0104541852176463,0.00033313477758834,-0.011052620909646,0.00895634037613346,0.00251395754562744,-0.0033198851063726,-0.0162723916354276,-0.00211095161698893,-0.00997862781066583
"2635",-0.000246946507627022,0.000226743735882273,-0.00147987635983204,0.00219630612481714,0.00204255262547104,-0.0000929136077107984,-0.00394764557882199,-0.00258485360419725,0.00287694195295307,-0.010799137029343
"2636",-0.000452798604804738,-0.000906550664983463,0.00203786751070578,0.00511314565961385,0.00219484122542357,0.000928730137329303,0.00198174857482747,-0.00414603915917855,0.00337496633584977,0.00145565913800816
"2637",0.00119422725604879,0.00340300837603924,-0.000739595308469787,0.00532946385358346,-0.000469384710851006,0.000278419537845354,0.00395545253556984,0.00442371498535832,0.00428861426654237,0.00436033063266361
"2638",0.000658106463446995,0.00339127329111566,-0.00277515856083066,0.00963860330116684,0.00375653077142335,0.000834799951527909,0.00640233589570038,-0.00207283226860033,-0.00895921460269622,0.00217088652750053
"2639",-0.00805625498013074,0.00247854770355893,-0.00241185774635211,-0.0116945671781526,-0.0106814685847428,-0.00491235087972963,-0.00591213103636745,-0.00519194447524407,0.00380193474314017,0.0115524115461247
"2640",0.00895038860576491,0.0074175000309622,0.00446335989229851,0.00772764660200442,-0.0033099207327616,-0.000931490823722236,0.00136569420831645,0.00104400458308174,0.000757545673891968,0.00642396808240298
"2641",-0.00878888277766632,-0.0111557491812805,-0.00999805134243037,-0.0127005622180066,-0.00838155485267744,-0.00372919015198181,-0.0109114021993393,-0.00469264608189479,-0.00487806551929248,0.00425518775965816
"2642",0.0018645644709594,0,0.00336637967379771,0.00461167059476519,-0.00231227620718,-0.00233957356847314,0,-0.00209554263299827,-0.00253552231237308,0.0204803110442378
"2643",0.00169566276299538,0.000451169342021274,-0.00484619307602763,0.00579843764276089,-0.00321957068656364,-0.00367317496057795,0.0106558496349711,-0.00892378669162797,-0.0163531693701027,0.0103806233302839
"2644",0.00231199084301403,0,0.000187215505753402,-0.00192169550406418,0.000240998531692682,0.000754485194369492,-0.0112876263351912,-0.00158893618094136,0.00370403148260934,-0.015068498558463
"2645",-0.00914448953539038,-0.00360852486771113,-0.00730345909690511,-0.0120337541608667,-0.00827367531089329,-0.00188430726938471,-0.0174380183888598,-0.00503982075981779,-0.000429076564428699,0.000695472358283933
"2646",0.00648517403635696,0.00203714481477402,-0.000565810604726713,0.00194884747945867,-0.00599372179926005,-0.00160468839538552,0.00485154240137176,-0.00106629860653629,-0.0102172404033893,-0.00972898790088284
"2647",0.00107382820780044,0.00225897595398572,-0.0026424040852695,0.0094821749011238,0.0014667458377966,0.0013237763325078,-0.00736970159406458,0.001868163413971,0.00164817836266629,0.00421046853524154
"2648",-0.000742656566059097,0.00135222438483185,0.0068129134632644,0.00818877291389941,0.00170857687455972,0.00132163649059924,-0.00115201602664039,-0.0061266845838821,0.00129905602061964,0.00978337842656662
"2649",0.00751479841871072,0.00855287671231553,0.00695479401550037,0.019350187457204,0.0069043883592117,0.00292329544632253,0.0125592570187354,0.0069684235707308,0.00354606460267948,-0.00484429563586741
"2650",0.00168024031774605,0.00423996933645299,-0.00130661196789217,0.00492161797262192,-0.00629247820739576,-0.00103428548709705,0.000379860484241767,0.00452510274548423,-0.00180986815314899,-0.000695400785539535
"2651",0.0046641056218899,0.00622230573685134,0.00242987082172164,0.012593256101108,0.0012178354694703,0.00141166027341155,0.0101213329676033,0.0135134078825567,0.00820235710585404,0.0111342268915033
"2652",-0.000122124473858842,-0.00154595701699711,-0.00130520848532278,-0.0046061951207832,0.00275694337842691,0.00122196760570681,0.00400819561686427,-0.00235307124192063,0.00445323296531375,-0.00344110942841314
"2653",0.000529469765998103,-0.000884883610975717,0.00522777406657493,0.00300786443131829,0.00873277745439571,0.00366060397680323,-0.00249519498592943,0.0094340229913521,0.00699121828807892,0.00414366093869045
"2654",0.00541397051634651,0.00199252008747086,0.00408619732501592,0.00830455444909739,0.000400753364200757,0,0.00800394853181219,0.00700961170151393,-0.000253992039166984,0.00894087224434292
"2655",0.000445328134861311,0.00552363757864138,0.00369956538323235,-0.00114401852348367,0.00288491791493439,0.000280590655457047,-0.00397029241867086,0.0043824169812281,0.00135497965184661,-0.00136337802319941
"2656",-0.000890195772498492,-0.00593259612023034,0.00184298376289238,-0.000687040818165063,0.00423432022684489,0.00177671751834363,0.00211780632052339,-0.000256510039579272,0.00862655630288489,-0.0136518315761254
"2657",-0.000243139546357463,-0.00309483718231918,-0.00202354508283809,0.00297952545029267,-0.00389849790901431,-0.000653192488661691,-0.00261036328794928,0.00025657585386174,0.000419218507140329,0.00207609617564697
"2658",0.00243094388509779,0.00221737917276554,-0.00350228380531203,-0.00251362868035343,-0.013019024103064,-0.00560376142183061,0.00124639486913725,-0.00154008591562893,-0.00326879562934856,0.0110497861959944
"2659",0.00004046750711173,0.00774339559958115,0.00332956250041172,0.00824738037952089,0.00161855450207127,0.00319308225889592,0.00535204271428324,0.00437014627097887,0.00807264561171617,0.00956278073642225
"2660",-0.000929670416769723,-0.00461030944993279,0.00331862877971778,-0.00545334299985967,-0.00492859196670126,-0.00159131081820518,0.000866537891226704,0.00179174842723406,-0.000750717402837386,0.0060892964033703
"2661",-0.00117310002483861,0.00110279713452899,0.00294003911957152,-0.00045694114894046,0.0059272334944287,0.00168767582148432,-0.00210274169306268,0.00383268824602245,0.00751315629423854,0.005379955507687
"2662",-0.000566933446813134,0.00264367474048122,0.00329797491808526,0.0011428750990119,0.00121057979145189,0.000281001925355628,-0.000123837579239283,0.00152670143586575,0.000497124857119502,0.00602005367344782
"2663",0.00222883082357828,0.00483422456970706,0.00584372181839021,0.00296805874005535,0.00702128828873994,0.0024839860623842,0.00446309038713433,0.00330385110791687,-0.000828140786749532,-0.011303174426881
"2664",0.000485153771637492,0.00109327485468547,-0.000544773836603452,0.000910432279300988,0.000561647096078977,-0.000935091037280622,-0.00629480549468087,-0.00253289250411703,-0.0020721093730276,0.00201745736003356
"2665",-0.00193987016425046,0.00152907250372425,0.00254317691005546,-0.00409361919403362,0.0103439580913995,0.00346282191866232,-0.00347767256331177,0.0012696472472209,0.00157802322960099,-0.0073824498756202
"2666",0.00182220842570979,0.00196296891110181,-0.000905963959782596,0.00365390834205082,-0.00849209429430131,-0.002704864448553,0.00336527856678992,-0.00202908023435067,-0.00779495838112476,0.00202830017005384
"2667",0.00185916275554532,0.00108837067232814,-0.00036268011231666,0.00682577784843352,0.00112067819332107,0.000561171531807014,0.000745249556049599,-0.00355781888778961,-0.00117007937868652,0.00202433339157682
"2668",-0.00246097211537388,-0.00652314776581264,-0.0010884729684264,0.000225992260157071,-0.00359809451811333,-0.000840988850449809,-0.00546163897741092,-0.00382548666041993,0.00292861680313594,0.000673322171594659
"2669",-0.0000404296961631356,-0.0013132520322876,-0.00617514530841046,-0.00903735857784704,0.00545668202083083,0.00121604447510504,-0.00174745097415496,0,0.0120974218913947,0.00672959153000807
"2670",-0.0141152448918367,-0.0149024915623966,-0.0104166062552177,-0.0237119124979532,0.00853952761753551,0.00373724244712492,-0.00762700883403933,-0.00972859536154702,0.00741901751576979,-0.015374396255745
"2671",0.00147671774441749,-0.00200217660450175,-0.00147741668438484,0.0023352693497698,0.000474645148789365,0.00111689297850881,-0.0047874723355178,0,0.00474594554247565,0.00339445675241579
"2672",0.00991315749221977,0.00735612993224066,0.00739782030394753,0.0102517679627521,-0.00514119277937974,-0.00241744954209122,0.015318197949183,0.00672182342423544,-0.00708529190418361,-0.00879568904694039
"2673",-0.000121574852535278,-0.00110645775601792,-0.00128509955099232,0.00115315458489529,-0.0042136276422593,-0.00298244852785856,-0.00286786002173778,-0.0048794234828835,-0.00770993286925747,-0.00477816212774163
"2674",0.00174442952614351,0.00531694187724674,0.00330873352210448,0.0103663142193597,0.0036726223456176,0.00186967425895634,0.00437677433548833,0.00851622646554606,0.00735658768333813,-0.00274344684758798
"2675",-0.0155909211398789,-0.0125605406702601,-0.0067790070293885,-0.0127680483545705,0.0074776137256658,0.00354562349220555,-0.00684781689225367,-0.00639715015232667,0.0050873470479853,0.00275099405355195
"2676",-0.00156316457462413,0.00066936559595776,0.00442728699882,0.00854507063859167,-0.000237016981737059,0.000186077088447645,-0.00739619228967958,0.00386316574434509,-0.0015511062380783,0.0178326868731391
"2677",0.000782738570780817,0.000892113592482202,-0.00220384791861916,0.00366387559399284,0.00244845537966243,0.000650706529586653,0.00896695602653041,-0.000256710063049503,0.0037612345765845,-0.0121294223954782
"2678",0.0104569944785529,0.0057930921149274,0.00202460472124288,0.0111795865948021,-0.00386069999049876,-0.00195091888672305,-0.000876096636783785,0.00179634612666213,-0.00448031110328595,0.00272854600406491
"2679",-0.00358520127092521,-0.000221498675187615,0.000367420217837644,0.00473819682208965,0.00680191905222749,0.00344396895794419,0.00826840867071454,-0.000768404752416796,0.00376400461307602,0.00884355670473025
"2680",-0.00233071954129804,-0.00132945275996066,-0.00514139955757087,0.00314397336631611,-0.0036920788067214,-0.00157673236051503,-0.000993995080555643,-0.00358891753256763,-0.00309771750383503,-0.00067436901525264
"2681",0.00233616448551621,0.00710010734645317,0.00332224588584795,0.00582040916624837,0.00386323090470952,0.00167196589442131,0.00472644085984908,-0.00128633623187835,0.00367975301594758,-0.00202419449601332
"2682",0.0000408113385552689,0.000220373144092623,0.0011037483717955,-0.00356093731937857,-0.000628219277000408,0.00092784776403243,-0.00507553991203691,0.00309118931269148,0.0158872741712119,0.000676053664256049
"2683",0.00114484051749297,-0.00396475647143568,-0.00202139079060126,-0.00178701026281025,0.00322235325235409,0.00231673461295245,-0.00149319718797536,-0.00205464342199746,-0.0021654021627171,0
"2684",0.00473750489782976,-0.00176930462831459,-0.000552420750399518,0.00156625109829589,-0.000313418757849404,-0.000832106484615736,0.00535845705281845,-0.00154380744156701,-0.000482213478254612,-0.00743240066882345
"2685",0.00601616830276219,0.00731078617567094,0.0079219264592747,0.00156399256353579,0.00297796846741316,0.0015731547520148,0.00644495055335215,0.0108247243898669,0.0117401012243479,0.0279101820157066
"2686",0.00141413337123031,0.00219905243840413,-0.00402106618215214,0.00736118616300607,-0.00764924735817385,-0.00294270956018849,0.000123232230007986,-0.00382463084077456,0.00190747099030353,0.00132448516535044
"2687",-0.0071822151617198,-0.0063636964782201,-0.00440453674104513,-0.0130648161361986,0.0158579587333882,0.00696012823325232,-0.00209314770381275,-0.00102360269523349,0.0111058307330769,0.00198403176737982
"2688",0.00341379757470439,0.00706698856664167,0.00423964013301248,0.00650674559192788,-0.00613539236209615,-0.00239595754130772,0.00197406266284617,0.00614884268760862,-0.00509964698807197,0.00990112731437764
"2689",-0.000121333496529985,0.0089912922443971,0.00587365977921239,0.00735616813996631,0.0102367531277343,0.004341638688385,0.00652742547551521,0.00814873306908925,0.01040932908145,-0.000653653071059468
"2690",-0.0011747321340706,0.000217403556616036,0.00310226013536963,-0.00663867043776079,-0.00216576415441316,-0.000735720568207032,-0.000611883028083349,0.000505420452520555,-0.00124876292637321,-0.0111183607233376
"2691",0.0106657895577305,0.00760530424850847,0.00454791071242133,0.0133660738347574,-0.0119381222887043,-0.00570705722103404,0.00844756599673957,-0.000252745761649575,-0.0139095021183909,0.00198403176737982
"2692",0.00337077427876387,0.00452875859730373,0.000724252617180454,-0.00109915992224308,-0.00525643300430856,-0.00240712903856388,-0.0100765205928909,-0.00429268900170843,0.00293205479147218,0.00264029608816352
"2693",0.000479920270305634,-0.00601115256179829,-0.00199043743718785,-0.00528153824431399,-0.00394346845744331,-0.00204123180125981,-0.00367908558394237,-0.0073548606863969,-0.00750629752696419,0.00460829992672163
"2694",-0.000319730117941619,0.00323984068423622,0.000181297698183647,0.00265471965681052,0.00411754034018408,0.00018581584336963,0.00615458728202123,0.00204390421318257,0.00437865612309007,0.000655366512221311
"2695",0.00134607497450356,0.000430596043653697,0.00145038363402228,0.00595765753177235,0.000393982280732397,0.00120886383723295,0.00415946009495416,0.00324036384996851,-0.0049936983197939,0.00458415661069123
"2696",0.00212686275945617,0.00193668671828173,0.000180926721635277,0.0035096434422246,-0.0057542849193184,-0.00390054826334274,-0.00536069832402941,-0.00281968994163939,-0.00932046530168462,-0.00130376311982083
"2697",0.00100113585005612,0.00472511299926537,0.00579189538606006,0.00218561644096082,-0.00245774612157357,-0.00111845919444864,-0.0077165668876461,-0.00308488402037255,0.00209072047209125,-0.00195826488688433
"2698",0.000360055839626172,-0.00299277192873426,0.000359873684092626,-0.00458008517888031,0.000715252710083103,-0.00195976357878613,-0.00246910901659481,-0.00257866660881534,-0.00802439396506838,0.00850230752397341
"2699",-0.00267937024950793,0.000857660845482888,-0.00395756201245245,0,-0.000555803850095238,-0.00130922254748556,-0.00321728517252551,-0.00698021921770875,-0.00760397166468274,-0.00389106408858941
"2700",0.000200585557960986,0.0021422573226173,0.00108376585898862,-0.00569677646657951,0.00286069127126787,0.00177908260918636,-0.00595904617893583,0.00442580913925994,0.0045647049233779,0.0039062636106455
"2701",-0.00204459109074562,-0.00769566323515347,0.00216480850546685,-0.0169678115838858,0.00625996847488541,0.00299106938150051,0.00537039275355533,-0.00544327248495557,0.0104673890046638,0.0168611887231829
"2702",0.000602535472371546,-0.00301591263000622,0,-0.00268990241360501,-0.0018113281371438,-0.000839025503149848,0.00027538152862161,-0.00208488560430409,-0.0111619690930858,-0.00892858080554015
"2703",0.00389432481438345,0.00172859523696456,0.00198014000568913,-0.00359634595531921,-0.0150675938374637,-0.00512950857878924,-0.00801603474341739,-0.00443992334568843,-0.00942013975491429,-0.00386108364400783
"2704",0.00119974053577998,0.00345122470334536,0.000718733637917746,-0.000676825436848105,-0.00296374451210391,-0.000187262136451705,0.00744968355138464,-0.000262239619274074,0.00188552217038396,0
"2705",0.00351518587949018,0.00752374686926305,0.000179451278659259,0.01151247600925,0.00224933692231155,-0.00121901996885709,0.0011279452822246,0.00708477303825483,-0.005155036454914,-0.00516788856168493
"2706",0.00433859848308327,-0.00192022717126594,0,0.00022314415014435,-0.00183113940497504,-0.00113782564355824,-0.00200292984174022,-0.00234495713987171,-0.00666232099584918,-0.00844151018349193
"2707",0.00214008965366586,0.00320648242649346,0.00592362169980376,0.0158410575511312,0.000965635416684263,0.00141198810781984,0.000752614647282268,0.00470090734544559,0.000496853535568054,0.000654869887072751
"2708",0.00118653669242463,-0.00170465343639781,0.0001783625295253,-0.000219568541018345,0.0000801727041708222,-0.000281999441705816,0.00639255000548711,-0.00519886202293063,0.00281383757653186,0.00130894998339981
"2709",0.00592513414254237,-0.0012806445795881,-0.000535197036823143,0.00746929128784579,-0.00377758806155337,-0.00103414101861021,0.00311370432270697,-0.0013064241283538,-0.0053643724579413,0.0111110931727056
"2710",-0.00113896511247391,-0.00085500292294205,-0.000535483626073141,-0.00501529585520832,-0.00282409967678976,-0.0012234489890488,-0.00360074613139894,-0.00183163634564298,0.00472949729661876,-0.0155139513659167
"2711",-0.00165100902889859,-0.00042774117279365,0.00125021201212938,-0.000657449123599219,0.00315554400961116,0.00113055974756704,0.00199379022622037,0.000262155574901612,0.00817578687507758,0.000656522276818006
"2712",0.00263826551010204,0.0106997799656545,0.00713514021220618,0.00986845878127807,0.00161342971540623,0.000376450817408891,0.00136778653627734,0.00707558202949476,0.00262123193608743,0.0118111334310549
"2713",0.00157094019304105,0.00254070440467302,0.0051364396301985,0.00456028557673838,0.00193241491302842,0.00112946284158277,0.00422274692782043,0.00572488508326163,0.00318626628780616,0.00194549867153038
"2714",-0.0014900898583472,-0.00190069352877853,-0.00123346911334854,-0.000432437999934199,0.00425981502623696,0.000939761035391173,0.00655452604809414,0.000517166387657753,0.00081438227205477,-0.00129448070386373
"2715",0.00121755394797396,0.00169284116070778,0.0123499612189721,0.00908309543224117,0.00720292152763147,0.00338040859364463,0.00221153001628749,0.00284463229670573,0.00756775170939661,0.00972125587305173
"2716",0.00133343600510161,-0.00253498176100242,0.00453122015507978,-0.000642867565873062,-0.000715056596732544,-0.00168447545298311,-0.00502618327902726,-0.00128939339917844,-0.00686479567113552,0.0025674912770961
"2717",0.000705105243962389,-0.00381201147642141,-0.0010409396666472,-0.00514700425751702,0.00127226315800377,-0.000375273363147355,0.000862435602853484,-0.00103279832687164,-0.00683096684694662,-0.00128045807361343
"2718",0.000978602718167521,0.00425188500683493,-0.00104187931328936,0.00237119188118551,-0.00659170006978038,-0.00253165992816828,-0.0011080435373656,0.00439390081643731,-0.00376647024727261,-0.000641082861988718
"2719",0.000273726427871379,-0.00169364851738529,-0.00226021329151105,-0.00881722796603135,0.00175896464559555,0.00103419222703405,-0.000739336120838319,-0.00128649917409351,0.00591765440811454,-0.00448993064839287
"2720",0.00516048224800825,-0.0029685665544138,0.00226533342823521,0.00368853998474616,-0.0106138633639259,-0.00413233678218206,-0.00320687675948261,-0.00438031418177498,-0.00637305340610395,0.0051545684159735
"2721",-0.00388938118639282,-0.00319004766593245,0.00243382316750651,-0.00799839558164739,0.00177458409200648,0.000942872098292469,-0.00470174783941568,-0.00879929212425501,0.00156238794866881,0
"2722",0.00175705764638168,-0.000640129090717756,0.00832464660729215,0,-0.00619953266638618,-0.00301484096983917,-0.00497281046064579,0.00156652965338111,-0.00385879300840419,0.0102564681117521
"2723",-0.00495014133093397,-0.00106738973649345,-0.00808399886624289,-0.0021789722318154,-0.00478018366592869,-0.0016065248374123,-0.00387284580844793,-0.00782061001711953,0.000164806722742883,0.00126895282363715
"2724",0.0012926915766216,-0.00235097738250478,0.00537538470984633,-0.00677014270075915,-0.00333779738855799,-0.00132497568392864,-0.00614577811312977,-0.00157656102733172,-0.00840540598937634,0.00443606490635928
"2725",0.00817620595210422,-0.0017138747520421,0.00758885418931698,0.0145117491637965,0.00661614985599956,0.00322224986430819,0.00454316593206583,0.00447368509817281,0.00473697324462785,0.00504724945748625
"2726",-0.0037251284529195,0.00579410551849846,-0.000342263778087104,-0.00628515641825811,0.00957471131776755,0.00359028565748765,0.00213556370729173,0.00104807291134179,0.00190235728862942,0.00251101593966951
"2727",0.0015577850186923,0.00512050667996933,0.00428079879334042,0.00937836942142067,0.000321621672320749,-0.000659068965524146,0.0018804668502892,0.00680448755237428,-0.00379756469406989,0.00250479097826695
"2728",0.00132227740572022,-0.000849104243377696,0.0056265404344451,0.00518593040109949,0.00445234182773979,0.000603692217812535,0.000750840351200655,-0.00441902817606388,0.00364633303466189,0.000624536740310377
"2729",0.000388420814954493,0.00254940917917112,0.00118683243441087,0.00128978808323366,0.00440892093887446,0.00132016560878268,0.00625146408676636,0.0039165979490845,0.000660564770369465,0.0062422403245177
"2730",0.0033387161328855,-0.00254292621972463,0.00237090410109864,-0.00515236920303475,0.00271372791077673,0.00160086901317613,-0.000621305916635895,0.0013005807761699,-0.00470335003377598,0.00620332494232834
"2731",0.00154766421174291,0.00212448487493355,-0.000168799818300647,0.011221374931971,0.00374062704410094,0.00122206975005779,0.011562916556578,0.000259409048572801,0.00853920555780463,0.0191123283471131
"2732",-0.000695346940217556,-0.00826791229300139,0.00794179266743211,-0.00640198939252756,0.00420270399441769,0.000375405960421737,0.00712872372984519,-0.00259659482527397,-0.00361695842799903,-0.00604964843524292
"2733",0.00170084349034316,0.000641177324395059,0.00620281919344245,0.00472493032316446,-0.00221092145452817,-0.00121997195495371,0.00671235202963771,0.00937250157281277,0.00346504416685955,-0.00182590324516907
"2734",-0.00362773091936797,-0.00704957631778391,-0.00833051165773502,-0.00619909987092115,-0.00284894079627374,-0.000375871759836444,-0.000363776645417757,-0.00232145852995636,0.00411082802213669,0.00182924326638534
"2735",-0.000309902728064859,-0.00150604410324462,-0.00739248422147565,-0.00430209055276021,-0.0150797118896748,-0.00507685425925586,0.000606374148621081,-0.00180973332506706,-0.00818799659841141,-0.00182590324516907
"2736",0.000929878440383947,-0.00452487778485189,-0.00440085365245357,-0.00216030466408501,0.00209531875751701,-0.000472591201482908,0.00363594768377284,-0.00492106925899716,0.00148601506198331,-0.00304873877730882
"2737",-0.00232257299626881,0.00216432874287342,-0.00527028932008733,-0.00671135309887894,0.00675469257619676,0.00141813562795479,-0.0015698882196814,0.000781061083902301,0.0020608359090073,-0.0134557875869372
"2738",-0.00500510953717204,-0.00453560562476585,-0.00734918920091643,-0.00523107286220958,0.010862741255184,0.00358725583097796,-0.00858726942314092,-0.00130042924984219,-0.00123390920095268,-0.00123984494504614
"2739",0.0085009708381929,0.00650911151876765,0.0154958059377404,0.0208150971089545,-0.00869160427237237,-0.00253975166885756,0.00670968213445122,0.00937482125059419,-0.0000823820086522931,-0.00310368377575998
"2740",-0.0029387602179457,-0.00129334331546327,-0.00491690757008123,0.00493659868213348,0.007412584374068,0.001320414639981,-0.00460476812697563,-0.000257909554525315,0.0120263507079679,0.0161893255167598
"2741",0.00170624750555315,0,0.00494120300855938,0.00512604967877905,-0.000395648258511239,-0.00160117059701936,-0.00206972483156742,0.00258054272708308,-0.0126160099901025,-0.0079657033931777
"2742",0.00654293725509825,0.00539588224975884,0.00915575160183879,0.0133871489294548,0.00316616184268415,0.000188917964616842,0.0071978300697455,0.00592027746394841,0.0016487017005804,0.0067942881877463
"2743",-0.000884576321978692,0.00364966779358311,0.000671999375899235,0.00251633513994087,0.00323501308259444,0.00320664286163841,-0.00278602657811355,0.0023029246361681,0.00921730706580015,0.00552146022906941
"2744",0.00230966138900235,0.00919794861258705,0.00822695931452633,-0.00209171234248029,-0.00275258310634041,-0.000846432502469963,0.00206505457729289,0.00459541546048792,-0.00252790514216528,0.00305072465542766
"2745",-0.000499244653825448,-0.00635864007889553,-0.00432962699266826,-0.0146719615148461,-0.00141965271733602,0.000658790710265977,-0.00412118854851173,-0.00101643663168338,0.00416940810987576,-0.0018248551037251
"2746",0.0101449343879656,0.00639933112224766,0.00301040246727946,0.00744536427329523,0.00134243380566135,0.000188234839759938,-0.00219080335081712,0.00432448073935898,-0.000162859233691082,-0.004265696046719
"2747",-0.000608667659080075,-0.00402716446741369,-0.00200092303428356,-0.01583623786513,-0.00985872254035347,-0.00319639317029585,-0.0012199550527211,-0.00658557029647444,-0.00626982340639715,-0.00673198010526599
"2748",0.00875493642933334,0.00106395962802708,0.0010024324930038,-0.010941892209768,-0.00334533929763459,-0.0031124795473858,0.0010991543161738,0.00484420354152015,-0.00770241717713527,-0.00431300522668032
"2749",-0.00207544790005698,-0.00361379574507503,-0.00450677732053417,-0.00563986297791874,0.0134943808159604,0.00369514212520738,0.00182999666139017,0,0.00404622632611429,0.00866337563776698
"2750",-0.00120995687754566,-0.00149360404960097,-0.0105633215462881,0.00196345140593968,0.000474106133216523,-0.000471876651379821,-0.00767193838341129,-0.003805960950367,-0.00337195504143284,-0.0122698975885782
"2751",-0.00359672804569233,-0.00363239660731685,0.00254189659012449,-0.000653270989964483,0.00497576790205989,0.000755573380545327,-0.00589006150596882,0.00382050163038317,-0.00709688067337855,0
"2752",0.000190123977521273,-0.00171571248115487,-0.00371867313053231,-0.0135075811856634,0.00345809403498687,0.00207631751459658,-0.000370315034806556,0.0017764186653435,-0.00207779255319152,-0.0167702126206949
"2753",0.00315290673924151,0.00257788818493476,0.00644719705161889,0.00287085745191384,-0.00783191712576581,-0.00178963913968189,0.00407508201073958,0.000759883712350362,-0.0131590072457732,0.00315851657128929
"2754",0.00545323914938423,0.00514254249910495,0.0047201021933565,0.0116714813340002,0.000078846082362638,-0.000754799254439775,0.00332065906549972,0.00379653363767729,-0.000084353111390878,0.0050378444325565
"2755",0.00301301850459157,0.0019185898783729,0.00335580261891066,0.00500665559058922,-0.00205231775755987,-0.000660765976932876,0.00110298260054997,-0.00176510290170606,-0.00396692258692799,0.00250629588749507
"2756",0.00176476413946669,0.000425465916426004,0.00183941102118457,-0.00671435223189976,-0.000395353248998642,-0.000850594391799797,0.0040406672471025,0.00303111920599974,0.00118634012056029,-0.00875007309041997
"2757",-0.000112335484871218,0.00212676683973667,0.00400613270487082,0.011993070450075,0.00751704438661216,0.00406651336555974,0.00207336519524493,0.00956941547733758,0.0086330595237738,-0.00441362391405054
"2758",-0.00408622995128016,-0.00594226374459028,-0.00465517803624971,-0.00732612172945091,0.00424102414655159,-0.000376946818622104,-0.000608514115397307,0.000249353298920507,-0.00201391293134034,0.003166583158283
"2759",0.00832748575963804,-0.00106738973649345,0.000501118606927919,0.00217071359304644,0.00375391021967997,-0.000188321796066537,0.00414015286418312,-0.000726835204406862,0.00210207685192976,0
"2760",0.00634112031443568,0.0132506551761458,0.0120200558964074,0.011262600189287,-0.00911595327942616,-0.0022615344821596,0.0055785074351169,0.00978429893774302,0.00461489343849641,0.00441919659547785
"2761",-0.00384043604492956,-0.00105464715164316,-0.0101459359118562,-0.00528343029170353,-0.0129736378901075,-0.00453325177686148,-0.0192564610113072,-0.00322994653453612,0.000751666230226267,0.00754251726589228
"2762",-0.000524128945376123,-0.00401185861603803,0.00134195712626428,0.00131145256333309,-0.0110730768282545,-0.00294156367187248,-0.0104387765562776,-0.00174472659348435,0.00267066432982821,0.0056144599261303
"2763",0.00205965743950154,0.00420375934602113,0.000670192274732306,0.0065488581569304,0.00582821605455242,0.000705206027636684,-0.00364179873667636,0.000749063388584714,0.00141500750303813,0.000620211184653829
"2764",-0.000261454147501228,0.000849928314172743,0.00468770042386457,0.00845802421419029,0.00136429080269274,0.000381277479735376,0.00630179278559129,-0.000498982528526204,0.00523650578067514,0.00433987205688369
"2765",-0.00119615340994172,0,0.000499959562221264,-0.000860230186418787,0.00296557462001612,0.00038067284694554,0.0048850155728013,0.00149769490917118,0.00686286577041728,0.0148148021084444
"2766",0.000486393093122039,0.00148620190855753,-0.00133248442615108,0.00258291245852194,0.0130255045890948,0.00428267664091031,0.00361434827349472,0.00648071022593255,0.00377766289999992,0.00243299406141095
"2767",0.00205754409837389,0.00233194272031767,-0.00233479041107731,0.00686984130997037,-0.000867777978241446,-0.00123187940547931,0.00583710230565138,0.00346689854913373,0.00507236345236772,0.00485430284159838
"2768",-0.00377050748960028,-0.000422941732748372,0.00183884562288483,0.00469086937655017,0.00157908708955201,0.0016127813579383,0.000247123697081131,-0.000740403489150387,0.0065120391780551,0.00301940706457482
"2769",0.00715738253031306,0.0067711028400963,0.00600693450716516,0.0188879207616086,-0.0107993961026042,-0.00331548660536662,-0.00506101901778311,0.00592733047153238,0.0121310147653697,0.00481637198410567
"2770",0.00632503446220034,0.00273221254936207,0.0137668161689519,0.00958144022710417,0.00478124389940815,0.00104530887563481,-0.0016129394166744,0.0056470652651488,-0.00263685173572759,0.00599165342118746
"2771",0.00421481850537941,0.0121567735683563,0.0122708915232557,0.0049514512350699,-0.000158556382210628,-0.000474431516878537,-0.0156581179565506,-0.00146475832944937,0.0051273754206056,-0.00119116894609306
"2772",0.00666397656209883,0.0068337265985785,0.00274782632482529,0.00862248144273225,-0.00285548117580137,-0.00123488450753972,0.0010099868784843,0.00440086268108519,-0.00103616292871167,-0.00357789130999808
"2773",0.00182886147543271,-0.00267376955682597,0.00580270346855039,0,-0.000636445059463364,-0.000475632592395248,0.00567543217355881,0.00024324867822223,-0.000159610625395157,-0.000598312713800175
"2774",0.00226336679492922,0.00144362073293092,0.000640936515176715,-0.00162836156945989,-0.0133723615207723,-0.00475719214452763,-0.011537507028303,0.00146026549491873,-0.00462848144008432,0.00658673582176394
"2775",-0.00153000124928793,-0.00329500427364937,0.00640618986660857,-0.00632012833265827,-0.00121029578893894,-0.000286795871739742,-0.0121798105095708,-0.00680439161360125,0.00240516309456029,0.00356925525226215
"2776",0.00729605680099188,0.00702486105650957,0.00668357020198562,0.00615517407671806,0.0041193368864838,0.000669191773427613,-0.00346784875949657,-0.00122348554525853,0.00327923700935173,-0.000592638145727076
"2777",0.00651912268915744,0.0133359767097359,0.00316159169770835,0.00958394549874164,0.00168932246079057,-0.000668744255273412,-0.00811932844398366,0.00710462496029596,0.012117322829762,0.00652416725529137
"2778",-0.00341821241350282,-0.000809832552305823,0,-0.00383744260310526,0.00417608930595836,0.000478039975319255,0.0027286298687017,0.00316226529577657,0.0016540564087435,-0.00471419813690632
"2779",0.00953134582401383,0.00445794798908183,0.00803665921042351,0.0131791905986414,-0.0013595659849257,-0.0021984484823675,0.0071270677976325,0.00703195828026848,-0.00809938677517319,0.00118411653188644
"2780",-0.00168053964775183,0.00100867924358861,-0.00844146655279188,0.00120061520482584,-0.00928962909673725,-0.00316124198923817,-0.00977857990394837,-0.00120406950429175,-0.00221973998905778,0
"2781",0.00454953377467793,0.00483683741280316,0.00630613761349541,0.00819503813308597,-0.00525413656418017,-0.00259461813079931,0.00649677446117058,0.00120552103540739,0.00444936433776144,-0.00177407408737407
"2782",0.0081310461966142,0.00681907301840434,0.00422992588608606,0.00574940251877343,0.000974933780819587,-0.000385338401330371,0.00813328754839393,0.00650118267641475,0.0018193640534625,0.00236963602636964
"2783",0.00212245923248311,0.00298795529780072,0.00608426347039104,0.00473101198627068,0.00430275964022209,0.00289174852923169,0.0138299991223381,0.00406727143556718,0.00497431496290068,0.00709240651970733
"2784",-0.000388264940292316,0.00317769428254255,0.000310146823091051,0.00843642148606816,-0.00541599945571591,-0.00192208881856515,-0.00353646153182241,0.00619493503468149,0.0121778992157284,0.0105631140112774
"2785",0.000423644462378192,-0.00395941969079128,-0.00480550393537027,-0.000583770075023082,0.00820868623036053,0.00221435441135598,-0.00190128888770846,-0.00331546073837441,-0.00667547144802505,-0.00580700294982217
"2786",0.0115776929215743,0.00795057205544625,0.00732086461518611,0.013821396488829,-0.00370797757315067,-0.00297821308927781,0.000380853467928599,0.00855312615335757,0.000781480028276382,0.00759347409706135
"2787",-0.00662973105278397,-0.00986001284778293,-0.00850468114742009,-0.0151690142502826,-0.00695846978288206,-0.00250562659737452,-0.0128220380948471,-0.0150764932424094,-0.00562199547627107,-0.0028985109481735
"2788",-0.0102569909779516,-0.0067715400852375,-0.0127885394460747,-0.0136479190705624,-0.00586651021285478,-0.00231865924227714,-0.00540122576608371,-0.00478352462145948,-0.00431876724489622,-0.00697676784298473
"2789",0.000496480804670574,-0.000200402693238066,-0.00568724902696516,0.00869727454485747,0.00590112924785458,0.000290418391898806,0.015774336331591,0.0108147879570832,0.00670346198651117,0.00117094409959151
"2790",-0.00113481274167104,0.00180507512613026,0.00492537471805199,-0.0135213467322498,-0.01449262553554,-0.00515845315853936,-0.01667508437995,-0.0116502577991716,0.00329028588656044,0.0099413840415421
"2791",-0.0217699850933832,-0.0248248640146986,-0.0147035225530051,-0.025625756448228,-0.00927940980906772,-0.00370382564606242,-0.0102266077893811,-0.0204473136180012,-0.0131178879376496,-0.0162129851678451
"2792",-0.0418228207759749,-0.0412646485192778,-0.0473363469251706,-0.0350662107814823,0.00944977506094724,0.00821750669792576,-0.0321736583204816,-0.0351177062264281,0.00253184589391431,-0.00941735710162106
"2793",0.0197025085561982,0.0220556884553873,0.0242547442562946,0.0325373398520228,-0.00621317004426369,-0.00436595928493511,0.00351362198130722,0.0132347561093435,-0.0104964249901067,-0.0059416896181449
"2794",-0.00542493167664382,-0.0121517686053776,-0.00888019677985896,-0.0315120224675709,-0.00950343092516348,-0.00292371253231449,-0.00390548332389862,-0.00979658862861632,-0.00470566289772678,-0.0113568727483593
"2795",-0.0375087769115374,-0.0250264282474072,-0.0296997128071651,-0.0346504016659065,-0.00109390836184331,0.000879484080493764,-0.029471194872281,-0.0228310147823705,0.00152257391199151,-0.0102780351854992
"2796",0.0150215325970893,0.00348048636594633,0.0100889805270943,0.0159773120668247,-0.00631870860555928,-0.00175796450834764,0.0207548956084842,0.00882663108864112,-0.00168031681036196,-0.0146611405460728
"2797",0.0146845377306144,0.0123564131397067,0.0194684686997029,0.0157259614243384,0.00440884287264764,-0.000293160064924303,0.00300221964580372,0.00823466587507804,0.00480889648494576,0.00619967137823907
"2798",0.00248724693176028,-0.00214140580614963,-0.0122883242708391,0.00763516238601647,0.00447400640767159,0.00166354463852625,0.00761908999044403,0.00306275655545196,0.00566322870710945,0.00184840363382421
"2799",0.0134963528248906,0.0199571101424367,0.0151311953525595,0.0250474007792596,-0.0110933265419273,-0.00605705697048697,-0.00486089323168037,0.00610704539066464,0.0170526171152821,0.0153751344041695
"2800",0.0127598496753714,0.00736380420763272,0.00480280521912535,0.0205338095279526,0.00339909537195959,0.000294697462944526,0.00990483838412803,0.00354055048221036,0.00116984328690162,0.00181718054121949
"2801",0.000293121677161112,0.00104428214044217,0.0153288605567954,-0.00321928800575311,0.00542074857671726,0.00235830504498047,0.00846437507289166,0.00579637895522045,-0.00327158423151652,0.00181375993405042
"2802",-0.00626116613595018,-0.0110577143035286,-0.00811691670498738,-0.0137262686143003,-0.00438052157113744,-0.0010784810420239,-0.0123900824718449,-0.00501128349812996,-0.0134417084514044,0.00301758450131029
"2803",-0.00497428281396828,-0.00443047604907354,-0.00998352771476296,-0.000818766045457164,-0.0122683596163247,-0.00294384852179341,-0.0165925028029354,-0.00805837249148422,-0.00459437586492994,-0.00120347674362009
"2804",0.00129614138550194,0.00508590529229291,0.00462882068819193,0.000614534655617449,0.00299827943729247,0.00137801912880797,0.00932794868409981,0.00279250749446525,0.00509310026760779,0.00903620732628263
"2805",0.0159392782162027,0.00674667593824418,0.0146452853615355,0.0178096988586951,0.00888169779343961,0.00383327984803739,0.0169884363529951,0.0151900746687539,-0.001266856660328,0.00656719708467035
"2806",0.0116123039425045,0.00649223009999766,0.0129745075444161,0.00925184583840655,0.00033879479790988,0.00117460631623079,0.00347441865536369,0.0107229749844366,0.00245757097239219,0.00533812706251435
"2807",-0.0124864478476135,-0.0158136912574516,-0.0136087683606799,-0.0290953901846861,-0.00143854290871248,-0.00312917870326579,-0.021041333266447,-0.0217119821603428,-0.0104389089072101,-0.0100296031652974
"2808",-0.0101302343828886,-0.0109935916610695,-0.00876475423862078,-0.0143677679064963,0.00635579074765835,0.00235413019093156,-0.00244862368704835,-0.0103407166584467,-0.00103889557353709,-0.0107270933030973
"2809",-0.0145405847037886,-0.0106883546840206,-0.0289832054392388,-0.00187414263185781,0.00682636314336205,0.00430390028966121,-0.0031366558084277,-0.0030580733526423,-0.00223999200000002,0.00180720426467462
"2810",0.00515494867019917,0.00108038528617782,0.0112984599482904,0.00417273741213275,-0.00812938373235716,-0.00370938399439791,-0.0017783227829905,0.00996914353631895,0.00537201727572145,0
"2811",0.0115577240441347,0.00669112296369434,0.0045023086523146,0.0014544198935158,-0.00270376781146175,-0.00127372640777546,0.0112374108440363,0.00202484254736901,-0.00167476674116562,0.00601333289763395
"2812",0.00253513197443422,0.00578909015645723,0.00614202784132534,0.00933608881385672,0.000931890362432242,-0.0000978940572974318,0.0063695900243832,0.000252608494514028,0.0107844623741811,0.00358632258656688
"2813",-0.000366284828552721,0.00255800625581015,-0.00841435346047192,0.00102774565307184,-0.00110023405292992,0,0.00511708895578655,0.00505071836936932,-0.00640162812298772,-0.0107207044128849
"2814",0.00483893439800043,0.00170119017867298,0.00615640422717045,0.000205320823285948,0.00576231985954023,0.00206030495061116,0.00509093658435211,0.00427121884352477,-0.00238627901379029,-0.00602051145286409
"2815",0.0174025087024243,0.00466991529880945,0.00248042124046899,0.0213507954181713,-0.00657191120474698,-0.00215407824583136,0.00626525760817698,0.00150106733769739,0.000956809136609893,0.00969115162118062
"2816",-0.00125514723505804,0.00169013696587705,0.000989857290128127,0.00241210281654824,0.00576707352845895,0.00235508825041419,0.00503351340077729,-0.00299772189119951,0,-0.001799615516479
"2817",-0.00646282997279957,-0.00864787870793438,-0.00164793134925645,-0.00902342991242167,0.00505953313593888,0.00166370514453984,0.00158170950972902,-0.00375868770689136,0.00191172533127504,-0.00300482847068939
"2818",-0.00513170001516194,0.00255319852837865,0.00429177951753479,0.00161872113413786,0.00880945823918955,0.00195465922141236,0.000789712202600157,0.00653927377422137,-0.000636047071363111,0
"2819",-0.0010895443330915,0,0.00197240228831741,-0.00363621525787683,0,-0.000390077423138901,-0.000262949374479016,-0.000749306505548053,-0.00636431996096221,-0.000602764527766642
"2820",0.00108447395590328,0.00190985836480961,-0.0044292073220864,-0.00223047805664389,-0.00357637157389745,-0.00117084194396777,0.00591889517132205,-0.00248812191490144,-0.00240195352438821,0.00361883050760348
"2821",-0.0135305278477929,-0.00635445773959964,-0.0169714525681043,-0.0107700805210251,-0.00317158007472806,-0.000976942374728673,-0.00928364085666133,0.00428303118543583,0.00216697435259983,-0.0066105484132043
"2822",0.0017009287659997,-0.00127908258954035,0.00569905548109495,0.0110929159903432,-0.00401897648170257,-0.00195572388818477,-0.000791905438251916,-0.000501645160609798,-0.00448470398451106,0.00665453856253961
"2823",-0.00191936231925338,0,0.00133330351270611,0.00589173898113371,0.00109281249121795,0.000685983476249596,-0.00766092978482036,0.00175721822769925,0.0174563996051227,0.0180288471202825
"2824",-0.0249971664197948,-0.0217715705593039,-0.00915454321140441,-0.0333265085420358,0.00990948102072053,0.00411189198036932,-0.00579782630002068,-0.0122777949169216,-0.00395319408713168,-0.00767416064361603
"2825",-0.0213145652216349,-0.0065459836358891,-0.0209977126262528,-0.0202675164362683,-0.000748521639368005,0.00136510620262653,-0.0159285801933505,-0.00659566903172992,0.0129385454928113,0.00892313813065582
"2826",0.0273590766028611,0.0197672540760314,0.0142415608252715,0.0324163483180913,-0.00382788351470631,-0.00272616469118503,0.0126199261906048,0.0114913958396738,0.0052503565139852,0.00058967534721921
"2827",-0.0170117681262981,-0.0105535830757678,0.00236843462170078,-0.0181781207626273,0.010692289983639,0.00566255356627887,0.00270939291735961,-0.00580652284350858,-0.00615841133581552,-0.00412480965262829
"2828",-0.00295495416899128,0.0065303796231162,0.0113079944740968,-0.00504944288558262,0.00264497181847934,-0.0001940675659442,0.019319054071635,0.00761785743864518,-0.013804965311867,-0.00414207687878376
"2829",0.0127777743169735,0.00843423854205994,0.0126835984613056,0.0209346046901102,0.00486366370796065,0.00203936895605183,0.000265141236337696,0.00856845468916001,0.000477197157149556,0.00891265673453767
"2830",-0.0215847403680856,-0.013939609407268,-0.0201054631628766,-0.0180198102730161,0.00197295148191778,0.0010191897607057,-0.0137802762479838,-0.00849566001129864,0.0116861514294764,-0.0135452839627221
"2831",0.0128170976624571,0.00587211742066818,0.0126135913798595,0.00991353945848639,-0.0077124079202251,-0.00320033739413661,0.00658325070466681,0.00579662900330402,-0.0075436035275247,0.00537306070353027
"2832",0.010699074012225,0.00410811772232011,0.00099644254870479,0.000417762201778915,-0.00206740992390786,-0.000583418172511951,0.0112120420273054,0.00927062649086952,0.00118760092190962,-0.00415671294288755
"2833",0.00789199761988102,0.00968994385817634,0.00497758012114691,0.00250510943547244,-0.00745696581918376,-0.00253114184316494,0.000924034777942451,-0.000993029353676289,-0.0051403243607826,0.00477048083169485
"2834",-0.0222859336453107,-0.00447859632884196,-0.0156843187168947,-0.0195750622325752,0.010935835438308,0.00439166872859298,-0.00896742678645668,-0.00422460570007643,0.0046899521934034,-0.00712168600849572
"2835",0.00492833013379546,0.00921174620786469,0.00888969489488134,0.00106201835209885,0.00165165272791445,0.000194355498507104,-0.00173013414883494,0.00698769265457733,0.00340217583196578,0.0125522520913601
"2836",0.0159003768931463,0.0123114222438756,0.00548623707248774,0.0195203932629966,-0.00181377027789942,-0.0017487074981164,-0.00386530938896523,0.00669156990068021,0.00236558113862162,0.0171191926377148
"2837",-0.00524201219142129,-0.00670987268459877,-0.00248007982592979,0.000416196649284384,0.00355138839282931,0.000973057049539872,0.00227469141289993,-0.00147717537198755,0.00778790101192817,0.00754505613080703
"2838",0.00822709973862379,0.00654422008126976,-0.00165761187242841,-0.000416023501696894,-0.0073245878270547,-0.00359682741615985,-0.00947924039004833,-0.000246664365603166,-0.0116306142250363,-0.00403226212851959
"2839",-0.00293333124398187,0.00167775277087068,0,-0.00998952921878815,0.00232138507769397,0.000877958440503201,0.00350436624078632,-0.000739805939448335,0.00655499905492807,0.000578361080894707
"2840",0.00822192989342341,0.000628281880856729,0.00282252601279298,0.0012612107313581,0.000330920402092261,-0.000487270309892485,0.00483552659632958,-0.000493360383622243,0.00141231858954072,-0.0034682796207488
"2841",0.0106983711717255,0.00732356264040845,0.0038079585382258,0.00209950994584007,0.00272855444831821,0.000584744756297884,0.012966182376577,0.00691347317695312,0.000940241344673742,0.000580157907066337
"2842",0.000740318944097318,0.00332377432130082,0.0067623723110668,0.00859002657175023,-0.0079987063572573,-0.00389853651612448,-0.00171529942451187,0.0029428160762861,0.0007827632093933,0.0185506490623992
"2843",-0.00554752861663865,-0.0043478545601614,-0.00376803216165789,-0.00581631830006712,-0.00814633335427051,-0.00274010765268928,-0.0142764650853223,-0.00537913503770282,-0.00195541653430453,-0.00398412652387103
"2844",-0.00847945773041014,-0.00270332573045351,-0.00197351159736281,-0.0125366749176077,-0.00720729005432996,-0.00333640986411732,-0.00858263835497841,-0.00147491161870306,-0.00760188883388535,-0.00171426242459438
"2845",-0.000150027783544338,-0.00125099056646294,-0.00131814502729155,-0.0080405679489719,0.000252959057891022,-0.000984776022207701,0.000676532005359887,-0.00664709043042877,-0.00797594585744166,-0.000572402055533772
"2846",-0.0134673027677412,-0.00501045235724606,-0.00362970466154733,-0.00469287042546063,-0.00455734678870912,-0.00118240649654566,0.00243312307028809,-0.00148708857616198,0.0048559145473035,-0.00515456898568611
"2847",0.00247155170344993,-0.00356701131508119,0.00314625122559131,-0.00771534359810444,-0.00669762055870515,-0.002170400685642,-0.00215746407532091,-0.00297826311036464,-0.00649607051027323,0.00172709207715172
"2848",0.0101658246257326,0.00568540698669628,0.00610755609287872,0.0144708468842485,0.00699882478836056,0.00286741118228639,0.012161994308387,0.00896179478322834,-0.00350851595539381,0.00517234311863457
"2849",0.000938854912306164,0.00125640766683621,-0.00278918374047554,0.00617408312813961,0.00771336540435641,0.00167629563887428,0.0129506019709753,0.00542824322067137,0.00424100980842601,-0.000571629824671294
"2850",-0.00769063445410367,-0.00460057962359028,-0.002303359303099,-0.0071941712984992,0.00176641048986914,0.00108248229025398,-0.00303142062034678,0.00147246295041192,-0.00725102788844623,0.00457659625192264
"2851",0.00177688863868752,-0.00546219613626742,-0.000824534834878099,-0.00490204690536844,-0.00360162468457936,-0.00156620975474142,0.00700667790336507,-0.0019605762998407,-0.0070631433361632,-0.00569480027258995
"2852",-0.00671744929481921,0.00042249561953267,-0.00594155324906209,-0.00792447880160541,-0.0010979007073566,0.000197303949205807,-0.00341327265367897,-0.00785663486117472,-0.000484981007881191,0
"2853",-0.00220365808776046,0.00358942628389314,0.000996128933526963,-0.00215888707950085,0.00448081292970381,0.00256499003999155,0.000395351056840187,0.00470185130204404,0.0050950019394258,0.00630014665445522
"2854",0.0129462183589597,0.00189356309769595,0.00729806023842317,0.00454354450430627,0.0015150761069338,0.0000980675264470321,0.0105343713498565,-0.00123151037188296,0.00209206631873249,0.00682990607890632
"2855",0.0033834251132121,0.000840000474134239,0.00115267907295102,-0.00581532986334188,-0.0015967959025418,-0.000491632248172835,0.0054731707670399,-0.000739805939448335,0.000240878430697755,-0.000565341543789177
"2856",0,-0.00125886498712691,0.00312496652650052,0.00563263581316242,-0.000925810333747612,-0.00167347523499273,-0.00492486164221162,0.000740353657481485,0.000160520189451674,0.00282807382389816
"2857",0.00966582924400927,0.00693271942051488,-0.00852590845900003,0.00193867226126043,-0.00598227721597822,-0.00226765023408781,0.0061214321977856,-0.00271266917955715,-0.00208679676015089,0.00902412904987493
"2858",0.0093505434865051,0.00479869110728837,0.00578796968773432,0.0208558047598593,0.00805256997254,0.00207517796703915,0.0091909712781697,0.00642953826034853,0.0068366282178618,0.00503079018948172
"2859",0.00305129290474215,0.00145340210156064,0.00756327330858619,-0.00168479461620408,0.0025223994625394,0.000098526275005506,-0.0041048115968163,0.00147407332809935,-0.00143792938169041,-0.00611782543922279
"2860",0.000476557412690148,0.000414787574506414,0.00554832719605325,0.00126571181804835,-0.00528395016398941,-0.00216919307390095,-0.00734149819921337,0.00318934618035494,-0.00408001599999996,0.0072746624522757
"2861",-0.00688702138405761,-0.00518148095950044,-0.0102240047666762,-0.0206489320005321,-0.0113828591665269,-0.0055342746267345,-0.0147918107333712,-0.0124726321560106,-0.0161458352662196,0.00111115316920229
"2862",0.00420499051534029,-0.00083328396554061,0.00295131851360142,0.0150602791200685,-0.0038380181620401,-0.00208673683694438,-0.00289724341162312,-0.00470514447922676,-0.0015512899685346,0.00554942804543024
"2863",-0.000844705093841935,0.00291912603025479,-0.000163481542810096,-0.0152607927168661,-0.00505114897624703,-0.00059748690125061,-0.00515134705393772,-0.00497640883204387,0.000572409840768451,0.00110373765033045
"2864",-0.00250008425739956,-0.00374224746389085,-0.0024526410570852,-0.00839421655004813,0.00860481939135727,0.00388572717629132,0.00225710056122885,-0.00300072072091795,0.000408654785807094,0.000551146903571942
"2865",0.00751846062546457,0.00605174980950562,0.00114750798826813,0.00607763164531283,0.000511967052256868,0.000694857425338036,0.0107298313573139,0.00652122607091576,0.000571840517217925,0.00771362090786609
"2866",-0.00278016481641663,0.000414849193183686,-0.00229224961897145,0.00345189758070674,-0.00153483837516033,-0.000396537685386056,0.00131071326637433,-0.00249198207239743,-0.000571513702526616,0.00109347875985599
"2867",0.00275135252761283,-0.0143063732230067,-0.00393819547255392,-0.000429909619510838,0.00725954282168995,0.00456418384042445,0.00850791740713652,0.00174879138923933,0.00106198019567105,0.00546159048228656
"2868",-0.00204865023839906,-0.00294482576542765,-0.00609548206418242,-0.00537739148905436,0.00796993476699059,0.00256812949983853,-0.00246604309147302,0.00174559465632607,0.00856858977828789,-0.00651827470529265
"2869",-0.00238264064779825,-0.00886088469226887,-0.00331515498710533,0.0041090000804036,0.00622490644633089,0.0039409046989638,0.00338272716912957,-0.000995748595916224,-0.00307465824337438,-0.0147621883463144
"2870",-0.0115009754479102,-0.0266069857372813,-0.00665227735747875,-0.0232609571246974,0.021902741815881,0.0107950278560258,0.00298229958451968,-0.00971850592121637,-0.00016230013929297,-0.0094340048311472
"2871",0.0133445380024191,0.0177126810783979,0.00703168953268207,0.00793821220651414,-0.00670811269369564,-0.00427197075263042,0.0126699859821062,0.0103172742859188,0.00146116565531007,0.0128852670219088
"2872",-0.00612582407709106,-0.00429742089527396,-0.00681633633891265,-0.000437502734392026,-0.00164728997686769,-0.000487303327743271,-0.00178743414771065,-0.00423430470448694,-0.00218857901786706,-0.00276550571138057
"2873",0.00981767644015252,0.00820034690831828,0.0068631176571976,0.0140075959969066,-0.00528369063506084,-0.00369467674921931,0.00345296868647549,-0.000250012028962132,-0.00495532095784434,-0.00665559702864238
"2874",0.00475146535119175,0.00256831771394261,0.00598496395432369,0.0101443832648258,-0.00723181850401544,-0.0035318721235682,0.00879436966338565,0.00850628569466516,-0.000979631006280179,-0.011725247698573
"2875",0.000727634728130866,-0.00170799988958792,-0.00181782583998613,-0.00769219656948505,0.00234448593269065,0.00255965443390704,-0.00126351761201804,-0.000992204471483182,0.00392248907601966,0.00169489199511852
"2876",0.0083605183248352,0.0100514597660437,0.00430462116181451,0.015073160601941,-0.00810299831755057,-0.00402626325230937,0.00113864371180283,0.00645622133105594,0.000569800579077073,0.00338416449252255
"2877",-0.000108031627448435,-0.00804575239772232,0,-0.0152735652070265,0.00968500103924907,0.00423995441733771,0.000631683287657614,-0.00764864242700525,-0.000488097957827893,0.00393474064972654
"2878",0.00295638255356745,0.00128072073713725,0.00296732272794431,-0.00193874021252616,-0.00300267540602828,-0.00137487501205857,0.00290432991689027,0.00198902164198689,0.00122090996890023,-0.000560017988806005
"2879",0.00132976907468252,0.0100191359509798,0.00312298023295465,0,-0.00184059184054242,-0.000983063920989902,0.00025188752790517,-0.0019850732882557,0.00178848058225367,-0.000560216466350849
"2880",0.00129267282105516,-0.00654283923743459,-0.00622639623611476,-0.0025902503771017,0.000251494814256015,-0.00059065616411158,0.00503532473783608,-0.00447534170592379,-0.00332713616829172,-0.000560415101785283
"2881",-0.00319103366167151,0.00212448257383535,0.000824347530323344,-0.00670846337066688,-0.000502661784625325,-0.00118131427427759,-0.0201654226171564,-0.00174812419838866,0.00301255495847585,0.00392579808687055
"2882",0.00251765620560507,-0.000635982325706164,-0.000988484255802557,-0.0067538624227701,0.00829968926096702,0.0031547376889971,0.00997059974830083,-0.00375287833153215,0.00154229236882375,-0.0111730327424138
"2883",-0.0012755976878861,-0.00615188463356386,-0.00527704688541009,-0.00789651522607793,0.000914433688753657,0.000786147953504512,0.00101256199750543,-0.000785632386428148,-0.0165342928319248,-0.0242939171124082
"2884",-0.00205690269238779,-0.0091783205456758,-0.00729431003484171,-0.0121600295916819,-0.000913598263723281,0.000491156883875243,-0.000885115806638304,-0.0053258979956593,-0.00189545910319633,0.00868564270287542
"2885",-0.0038327222031892,-0.00844301625929922,-0.0106025435886629,-0.0110384897774766,0.00582020470925837,0.00264996951625762,-0.00012653394337292,-0.00535444420442532,-0.0025596399755623,-0.0103329868542164
"2886",0.00170589421074996,-0.000222243720307547,0.000340194235066926,0.00432798546286106,-0.00876253204995425,-0.00323042829905784,0.00974561835320165,0.00281982411146031,-0.00447020684262733,-0.00116019641551013
"2887",-0.00626868338162212,-0.00778289768124085,-0.00374096895489739,-0.0140620047128914,0.00525391004070652,0.00265169470047044,0.00513919414518194,-0.00460115534591798,-0.0017462081864924,-0.0075492592332711
"2888",0.00182320713644324,0.0136708385401572,0.00494971684439172,0.0103518570197556,-0.0000830599781372898,0.000195956295543809,0.0063597421221504,0.00950165877963083,0.00241560177220479,0.0198948260359761
"2889",-0.0136130055342731,-0.0148129732975072,-0.013586917624913,-0.0134334187857085,0.00224027433326168,0.00137098748987663,-0.00346936622146377,-0.00661415529886733,-0.00373938021403952,-0.0114746066791805
"2890",0.00221409944100115,-0.000224431859121799,0.00585385834586627,-0.00392351231522559,0.00140727643144167,0.000488976735951496,0.00395501679792876,0.00409740395509517,-0.00525479193639833,0.00986655672432346
"2891",-0.00828436426975721,-0.00965215228217298,-0.00667574159840878,-0.0192307631799801,0.0094238293109723,0.00381243499550554,-0.00537789701063229,-0.0119866004336716,-0.00570182784333684,0.00517234311863457
"2892",0.00571747152801327,0.00249325309116055,0.00120622953537253,0.0085046360443537,0.000245864907873594,-0.00097399597107739,0.0106878287538643,0.00309752501272986,-0.0030359334957677,-0.000571629824671294
"2893",0.00143987945883706,0.0108522814175827,-0.00327012986893371,0.014991901655999,-0.00343896138888478,-0.000779711192177124,0.00248830299774316,0.00720513211443086,0.00363729484319664,0.011441608389076
"2894",0.0021379551666536,-0.00715719027888451,-0.0158867186716306,-0.00992399385231391,-0.000782252954780627,-0.000684208500468353,-0.00595684661890472,-0.0071535895565833,-0.0100295236404632,-0.020927723011414
"2895",-0.00353140335967317,0.00585717731587532,-0.0012283139585213,0.000699351833970407,0.00535634677634489,0.00254280167308041,0.00749051389684507,0.00591863897772726,0.0101311340893167,-0.00115526692314427
"2896",0.00815785149866466,0.0132139276411276,-0.00158119526929035,-0.00256244119364391,0.00286897348636428,0.0000978666250106563,0.0130112063269479,0.00690723439887408,0.0033712683797511,0.00578367033561245
"2897",0.0084583097838582,0.00486280262766225,0.00651069783435787,0.0137786815979142,0.00326921925795309,0.00087764622611064,0.00415885206830624,0.00685961950134306,-0.00159598484008439,0.00460028213185626
"2898",0.0090045860620962,0.0063793741323166,0.0138111934818705,0.0179682246578181,-0.00643574379902079,-0.00253388018205891,-0.008892482425915,0.00454217373504529,0.00243985358876109,0.00515173632649257
"2899",0.00359817057287226,0.00240433131790208,-0.00379381451787619,-0.00226293964438407,-0.0000821040288733199,-0.000781632112785591,0.00307291987280256,-0.00276327284179345,-0.00184642884017738,-0.00227787321992068
"2900",-0.00731433327573117,-0.0183165532169245,-0.013847978993315,-0.0195055058245853,0.00385408551050692,0.00205332460049434,-0.00306350596444394,-0.0130982441432218,-0.0108467249642648,-0.0348174624831071
"2901",0.00906608206011739,0.00888485406674011,0.00105316887974105,0.0136479036866912,-0.0000816677845814073,-0.000390021576353372,0.00294983028404894,0.00535988166523826,0.00416523294938154,0.00532240485517366
"2902",0.000787339819464661,0.00286218790593917,0.00929340896055453,0.000684573568380253,0.00253252981113339,0.00165928697565176,-0.00343128623195621,0.000507812557802412,-0.00440189632782273,0.00176480282097224
"2903",-0.000894104504672755,0.000439016598250186,0.000347481730034183,-0.00547312785178355,-0.00415578382509574,-0.00165653830322066,-0.0045500196565047,-0.000507554815093569,-0.00051014369092639,-0.0211392979429703
"2904",0.00404517332898702,-0.00175534146653578,0.0088571343194126,0.00733779152586345,-0.00188213251139635,-0.00058602043124989,-0.00531193120698015,0.000253906278901095,-0.0108039469807585,0.00119974367765274
"2905",0.00210373620119908,0.00241798164218276,-0.00154927736587518,-0.00113822576932954,-0.00401694267418162,-0.000781403134530789,-0.00471931093716449,-0.000761409451884965,0.000257989338303899,0.00898741846514817
"2906",-0.00377146768028602,-0.00350882950969988,0.000172387353531755,-0.0123063082622605,0.00633810107227628,0.00273721709542896,0.0101073089762262,-0.00558816592267031,-0.00429885657809059,-0.00118763226939633
"2907",-0.00114291352910001,0.00572192521330295,0.00310298746917725,0.0143055166666228,-0.0122690533516375,-0.00350955387547769,-0.00840021890143283,0.0109835584233924,0.00647612479882786,0.00713438888152895
"2908",0.001859388730995,-0.00262579524367568,0.00498359939304716,-0.00659697637731194,-0.0123387314778158,-0.00489113184351941,-0.00249162046936224,-0.00480045447351563,-0.00480437551139967,0.00354192497063477
"2909",0.00503206561333225,0.00680105438023548,0.00410402422008316,0.0146553970809096,0.0034377303048545,0.000687856452955771,-0.00487080071792245,0.00330052049481511,0.000344836206896515,0.00529404521019172
"2910",0.00852250854334624,0.00740909862630712,0.00647136094667911,0.0162490921267611,-0.00158756995210774,-0.000687383631689076,0.00815774475971187,0.00607266322060918,0.00551533087284284,0.0134581601662647
"2911",-0.00235926563223698,-0.00605654763412311,0.00253808233543062,-0.0111037245934639,-0.00192484553048977,-0.00108163873910916,0.00273880516272507,-0.008299756116946,-0.00779913438464175,0
"2912",-0.00677608695783272,0.00195858074650701,0.00303797771750203,0.00359309604217528,0.0016769926384832,0.00157465924445432,-0.00968356259090042,0.00152177623767669,0.000518312184114356,-0.00404145601756001
"2913",-0.00522350801642213,0.00260640409212165,-0.00757198419526428,-0.00156630471810926,-0.00343213126240471,-0.00127763179581641,0.00137881038750098,0.00177281406304353,-0.001554001527169,0.0057971412257396
"2914",0.00492931302969546,0.00411597121832408,-0.00762968680031517,0.0053788429181918,0.00545989938632019,0.0013775008855772,0.0171508537994756,0.00454974718346346,0.002939870247473,-0.00576372808007275
"2915",-0.00167065359042684,-0.00755106247583337,0.00649235099316736,-0.00891672968623669,-0.00814676965618133,-0.00236255594609569,0.00332311066590041,-0.00603924735727024,-0.00732820945474966,-0.0144927933996526
"2916",0.00544771721210768,-0.0091304033433266,-0.0056016578773358,-0.0132703313464081,0.00143507553798394,0.00118399876339614,-0.00331210417718264,-0.00278484388017475,-0.00538476641814112,0.00588239354001052
"2917",0.0042846226454929,0.00197445693757392,-0.000170750808167863,0.00775026933724754,0.00497349589928842,0.00256278179931946,0.0118152700642558,0.00406203622970724,0.00349284850225762,0.00350872377936784
"2918",0.00366726241336424,-0.00459826872031011,-0.00751231566041777,-0.00769066461509815,0.000587183962076798,0.000491512732538002,-0.00060813179057817,-0.00455124540560403,-0.00513397154775463,0.00174822784108608
"2919",0.00330223362003101,0.00791915753652983,0.00842932844193856,0.0102575434371421,-0.00519732034868403,-0.00206346958929993,-0.00352960960083082,0.00330199380369978,0.00227406625952842,0.00756249299486456
"2920",-0.000420189733206455,-0.00174585481003298,-0.00102352492264934,-0.00135379536807212,0.00101114602755725,0.000886383952740211,-0.00598521918845685,-0.00075948183368868,0.00279263470783264,-0.0121246057469363
"2921",-0.00136594491167241,-0.00349808934594753,-0.00375686944404663,-0.00293705805499078,0.00841807314354592,0.00275428881569728,0.00122896748493506,-0.0035470196108216,-0.00147947083876176,-0.00409111864171874
"2922",-0.00670015479271246,-0.0223782137557023,-0.0143983515651468,-0.0213008219146434,0.007262764313404,0.00431675889426142,-0.00895924873871856,-0.0142384086234916,-0.000435732969073177,0
"2923",-0.00374349716445244,-0.00269313559661877,-0.00591303161338774,-0.0164388788545115,-0.00207208779623835,-0.000293099874108416,-0.000495304212960734,-0.0046428986549506,-0.0150841657496876,-0.00528167780563416
"2924",0.00638061162235481,-0.00180009255852376,0.00402373390710764,0.00612054807698414,-0.00224221156256788,-0.000976999270339896,0.00545150534178029,-0.00259122569174774,0.000973804895306296,0.00176976566726261
"2925",-0.00746726123446617,-0.0171326916457107,-0.0121972061268161,-0.0287787587415663,0.00582653721022686,0.00244515528864531,0.00751701567748864,-0.00545599598360869,-0.0166268506235074,-0.0217903474683254
"2926",0.00809139964682037,0.0071102927387634,0.00546835125206191,0.00626354753842007,-0.0000827490343077164,-0.000292756693700547,0.00807239755260891,0.00705330082506395,-0.000809461267929579,0.00782656574689478
"2927",0.00352013853649757,0.00592110946999935,0.00333332767644468,0.0105339126053279,0.00124147597410262,0.000390473415075476,0.00897838231802006,0.00648487427933175,0.00927091825870252,0.00418166710267975
"2928",0.00214004160279169,0.00701834738735463,0.00402169519788687,0.00450134324093443,0.00669532759593139,0.00312193143367412,0.00156317397118722,0.00670121236917587,0.00499424788176883,0.00178462762613107
"2929",0.00234544406400117,0.0107913801206971,-0.000174200325966156,0.0127357691723415,-0.00336657905451831,-0.00136170563578397,-0.00672332727117597,0.00179200872078744,0.00292834319055202,0.00178144840409455
"2930",-0.000593680568823474,0.00333624944292832,0.00418051452505774,0.00791805269647239,0.00395455751879048,0.00185039911370155,-0.00556042269910062,0.00178903682857867,0.00221199793519733,0.0142265489565536
"2931",-0.00132798928026123,-0.00753720921266809,-0.00416311058080521,-0.0161735909090701,0.00155933631127025,-0.0000969398199147653,-0.00218806873055821,-0.00612255744874024,-0.00944645562231283,-0.00175333656073662
"2932",0.00601834394978318,0.00826451794918714,0.00348373521676471,0.0185532006761251,0.00196616829961904,0.00029139140786838,0.0051165561152382,0.00487673086191731,0.0174688685597737,0.00761113664734459
"2933",0.00789540141932288,0.0132921532078663,0.0151015335874842,0.0142956204977316,-0.00572383675109278,-0.00223531299661872,-0.0018180439515012,0.00791861762006274,0.00376657309857831,0.00348629761126173
"2934",0.000483246603521392,-0.00174918119620882,-0.00307792578083277,-0.00363720253512789,-0.00600389699586479,-0.00224033090397924,0.0106848899879575,0.00126681559475816,-0.00794132150942739,-0.00405309730294123
"2935",0.00538081207531826,0.00459918468149234,0.00360207070524399,0.00616004211989729,0.00132376537714918,-0.000292928162657025,-0.000961077615621031,0.00556824959476243,0.00457421710063333,0.0110464194354272
"2936",-0.00404832722084658,-0.00981027971412185,-0.00700745274503134,-0.0260770231136993,0.00214854997330249,0.00185538779748295,-0.00348725469962963,-0.0113264501078533,-0.00490366037400147,-0.00172510579944607
"2937",0.0000342921958782494,-0.0112285921364474,0.00206551297911783,0.00512225272299816,-0.00230884122991648,0.000194953975263479,0.00374087062661133,-0.00152747116060947,-0.00114393700408255,0.0011520579548232
"2938",-0.00172217756644932,-0.00823866165796805,-0.0123669316059342,-0.0194579991046908,-0.00578144614873255,-0.00228500876400173,-0.0105795551683415,-0.0114736466563375,-0.00510969949590867,-0.00575372044135014
"2939",-0.00269153808633327,-0.00583745204379282,-0.010608661732083,-0.0144105592641929,-0.0026661228966427,-0.0000979543535343241,0.0046172405639755,-0.00438504991408639,0.00345346674931357,-0.00405098955429095
"2940",-0.00300988074651243,-0.0049683942490315,0.00228510482726429,0.000958776059713395,0.00367560402693212,0.00205564427207605,0.00387050214429951,-0.00103605603502188,0.00194141369572898,-0.00581049601876982
"2941",-0.0019432961017477,-0.00817059828053601,-0.00613823028804095,-0.00502877788020129,-0.00848932940112834,-0.00449349247596098,-0.0121686853234357,-0.00674271204010124,-0.00273029766839628,0.00233778208098223
"2942",0.00173829324813402,0.00892447655316331,0.00229397598097636,-0.00986761331554453,0.00369330710218585,0.000588819863478918,0.0063421150097196,0.00104429046660615,-0.000706535351765347,0.00349849440394534
"2943",0.00329745983131424,0.000453577826141416,0.00211269635556022,0.0021877102578749,-0.00761054329323263,-0.00362853046001443,-0.00206050968612004,0.00365156142570622,0.000618638963877371,0.00987802264203652
"2944",0.000242287270365127,0.00385398211431975,0.00193252981082548,0.00509324388332266,0.00235964982444292,0.00118108024794705,0.000850330865219462,0.00545726555242099,0.00839071711366635,0.00690439346752192
"2945",0.0059143718472241,0.00722678732238702,0.00771524546000113,0.0135136368270001,0.00151340848029169,-0.0000983775318521563,0.00594591010963375,0.00361864692286384,-0.00359110105266014,-0.0108571717928199
"2946",0.000172017367982225,-0.00224218924851982,0.0113101975962075,-0.000952384197535516,-0.00478523126683572,-0.00186787322186399,-0.00808220538860782,-0.00309034569541267,-0.00650496648198018,-0.00635450319835917
"2947",-0.005294282314943,0.00269669693858243,0.00051623595361372,-0.0090562500343867,0,0.000196928838708699,0.00352669504911596,0.00258342874332707,0.00522035051903247,-0.00116289437072703
"2948",0.00542622645662494,0.00515457196554658,0.0239036946898419,0.00962001736592022,-0.0104597304958937,-0.00413629980217434,-0.0035143011805413,0.00669901192334899,-0.00149633833732643,0.00931320734642194
"2949",0.00106550651783466,0.00222969106137638,0.00352703553878886,0.0138161251222619,-0.00596691062358878,-0.00168137023138315,-0.0132554148649023,-0.00358310040304266,0.00387865825319711,0.0063436269774495
"2950",0.00810399422485042,0.0180199821257478,0.00267782696580698,0.0110431968543943,0.00463067693190178,0.0000990562501268499,0.00998283371978581,0.00796280702092278,0.00342465762446409,0
"2951",-0.000913717598463371,0.00043702463620332,0.00216991514095666,0.00464793596539637,-0.000426765938975282,0.000396267663162142,-0.000488141840056966,-0.00789990162876852,-0.00682592999455489,0.00229223237918608
"2952",-0.0033220462536433,-0.00480551203005752,-0.00449698083657923,-0.0113346873852362,-0.00256189272427065,-0.00108908949600484,-0.0175802927846511,-0.00363370940916852,-0.000176200549408811,0.0148657296621684
"2953",-0.000927764736132763,0.00570676254228153,0.00752891112892518,0.00397740537521996,-0.00102754020838969,-0.000990997825952133,-0.00161562603081511,0.000520960813086502,0.00158633117488027,0.00225360625707682
"2954",-0.00299222803177124,-0.00152768542268467,0.00481553512866739,0.00209744488717556,0.00702793022941473,0.00327406506122863,-0.00915052348452927,0.00364497412513654,-0.00527935758417319,-0.00449707787132436
"2955",0.00279423985136429,-0.0028416106876884,-0.00264417689167384,0.00488368930950589,0.000680895730093667,0,0.00266401583847697,-0.00181598563830876,-0.00884564328582993,0.0045173929391471
"2956",0.000103030976852603,-0.0120560973157002,-0.00198836900983113,-0.00671145709727794,-0.00263648918652459,0.000494223610771449,0.0123985651939502,-0.00597714038859021,0.00633644784462883,0.0101179045278676
"2957",0.00347443016658056,-0.000443784543227688,0.00680727158259242,0.000233114132708545,-0.00734145186627433,-0.0025354302660533,-0.0082477066821095,-0.00261413121893039,-0.0016850123858636,0.018920451388869
"2958",-0.000582891580144684,-0.00532729375464069,-0.00230876034615191,-0.0125786351757077,0.00611267688335393,0.00258180275453901,-0.0013860495101583,-0.00996081986790243,0.0115483965532557,0.0032769655314917
"2959",0.000548916107523612,0.00379361414247392,-0.00876031430284863,-0.00825661886464868,-0.0173710992056993,-0.00742794044161532,-0.00694007819726294,-0.00529527424288656,-0.00395191875071776,0.00925425988695894
"2960",-0.00781595122312118,-0.0131168220587201,-0.0135066901799198,-0.0249761987618015,-0.0070539824302267,-0.0025942710538065,-0.0100380932468805,-0.0188979565084041,0.000529051323030272,-0.0107876155675189
"2961",-0.00559697247011559,-0.00698356388127841,0.000169007203053573,-0.00365949250137498,-0.00859496595097164,-0.00240103807520331,-0.00128372221395012,-0.00189900160486223,0.00281988008054612,-0.00218110757682066
"2962",0,-0.00930131679799473,0.00439412303544495,0.00146915296724637,-0.00336145051158565,0.000401255121219135,0.0132375088672902,0.00462073226467918,-0.0110720735218258,-0.00273220340393854
"2963",-0.00145915237982241,-0.00114495769254785,-0.00572107396498189,-0.00366754538905723,0.0101188051200378,0.00190448384888109,0.00215624598561837,0.00865793340554566,0.000533117109177805,0.00712324725195068
"2964",-0.0316631407588487,-0.0194863534993317,-0.0245387517141701,-0.0296931507380268,-0.00272425231090934,0.000500177309976868,-0.0150613257568177,-0.0179718969360335,0.00248666967116651,-0.0195864096426023
"2965",-0.0220266277207172,-0.0126258055047875,-0.0180430430716371,-0.0101163459436877,0.0121599159284445,0.0040999873909231,-0.0272424388095432,-0.00409737688968093,0.0256910176920009,-0.0149833186461571
"2966",0.0138883899050801,0.00189456695698653,0.00229674022630433,0.029381700311466,-0.00348219356459534,-0.0011948563745694,-0.00198144623390062,-0.00192005260700301,-0.00475035416091174,0.00788721601174891
"2967",-0.00561702622511007,0.00165442067713695,-0.00299660863246398,-0.0106726859329337,-0.000436889057888523,0.000598070879916035,0.00542680567093679,-0.00109909265718822,0.00668226138985695,0.00223597067338011
"2968",0.0218659365199874,0.01604517349859,0.0185643480590378,0.0250879471836001,0.00227254636757435,-0.0000997662457843385,0.0217219944854814,0.0198073651555934,-0.0017241120689655,0.00446184972113572
"2969",0.000178288329387932,-0.00952154904876357,-0.000694288889770078,-0.0122370241891204,-0.00592971391338404,-0.00288986008045744,-0.00489631225917786,0.0016186561757574,-0.0000863730547572272,-0.0088840601011867
"2970",-0.0144410815423558,-0.0164126865136246,-0.0180649823128983,-0.0262635890306195,-0.000350886828124675,0.00179889808483336,-0.00116527170515723,-0.00430911601279171,0.00112269625077555,-0.0112045023045214
"2971",-0.000542709888583959,0.00786647578168509,0.0021227870212448,0.00941473739094789,-0.00219366706476809,-0.00119708446173461,0.00764852382143499,0.00405711127142139,0.000776432035480168,0.00566582033804575
"2972",-0.00448881225723385,-0.00591292319831371,-0.00617832109645589,0.0108393836521843,-0.00131942720455969,0.000199691371261634,-0.0131226152296577,-0.00484897085754077,-0.00258600978215662,0.00112674514453537
"2973",-0.00509054122005692,-0.00713775220408586,-0.0115452409161565,-0.0109724766302115,0.00317025451091668,0.00259660280486917,0.00638778636202653,-0.00379002295411734,0.00587676091847511,-0.0219470914597191
"2974",-0.0302986927454122,-0.0282769595835076,-0.0319856924745601,-0.0322743888021586,0.0075491834278989,0.00537880806447677,0.00725396899155872,-0.0138586167202779,0.00231982990222379,-0.00690445268593698
"2975",0.0179405278977338,0.0128235763053226,0.0148506007417497,0.0192808060151362,-0.00418177568321099,-0.00237779962646001,0.0123455245581017,0.00909350465734149,-0.0022287158502069,0.00405556430793319
"2976",-0.017587293358195,-0.00413917782058759,-0.0128040537354562,-0.0115030546247896,0.00603659359047559,0.00446936311065982,-0.0235008294526332,0.00191144713493596,0.00317865114813309,0.0075013995081854
"2977",-0.0055402632538406,0.000244439161749099,-0.00926439600485041,-0.0173260453693882,-0.00226093931036642,-0.00009882377069792,0.0115779496311679,-0.00327074852481657,-0.003939359525718,-0.0103091969184586
"2978",0.0148185245100145,0.00855536600843476,0.0157097395019186,0.0194738066409266,-0.00496815082534374,-0.00217558230386572,0.0150463056428169,0.00464877824041676,-0.00438479072108655,-0.0052083811063095
"2979",0.0106808858001062,0.00799812935216959,0.00975869724266243,0.0108413280188648,-0.00508064605010305,-0.00247732974372872,-0.0103889358903267,-0.00816566586652534,-0.00561313456960799,-0.0133799887343048
"2980",0.010641830639275,0.0158692085988228,-0.00237052556661188,0.035750918647101,0.000926749541885874,0.000856003158337781,0.00371271872234713,0.0148188658017814,0.0128527570498871,-0.00707537594761776
"2981",-0.00592283800017002,0,0.00566631192418332,0.00641017501899466,-0.0124328532385911,-0.00557048934708493,-0.00854585254899032,-0.00459708411791271,0.000171525340946443,-0.00237526453879289
"2982",0.00551680141163535,0.000709935293166764,-0.00363513885639388,0.002694817962686,0.00392862136430172,0.000600273384538941,0.014665934269064,-0.00135825922307065,-0.00240033429232178,-0.000595229963322619
"2983",0.00632786639337057,0.00165559486421696,0.0113097718436566,-0.00171019175157183,-0.000622579881949026,-0.00109970893653233,0.00431095836674134,0.00788911677167969,-0.00283579953160262,-0.00416921391002356
"2984",0.0214089328648526,0.0129870921385065,0.0104617527745046,0.0188447201796276,0.00133487962888901,0,0.0126246849933245,0.0156546094178613,-0.0000861944149759264,-0.00239218884047798
"2985",-0.00181504223252626,-0.0114219413258506,-0.00642622794948,-0.0259428944320121,-0.0000887521516336198,-0.00140108801950556,0.000373936342836778,-0.00876992532914433,-0.00215461520429727,-0.00599530645430091
"2986",-0.00976814978720086,-0.00377258541306236,-0.0100611321817843,-0.018495646572353,0.00746592402670365,0.00390848938862276,0.00137104467876914,-0.00482569251705001,-0.0112281569461752,-0.0108564294470516
"2987",-0.0186852648009936,-0.0201182901969638,-0.0136115641135693,-0.0140702958894899,0.00652843521319268,0.00299501477247754,-0.00112012831466857,-0.00592654025201023,-0.00716281427770404,-0.00243899102184708
"2988",-0.00187113088627144,0.00748773044522344,-0.0036798753979963,0.0114678760482385,-0.000613784218886693,0.000796213999512352,0.000872157396843765,0.00785893919310809,0.000351865199652801,-0.0275061756106754
"2989",-0.00683674063957396,0.00119876057708068,0.00350882300752553,0.00604685771899161,0.000614161181327733,0.00208853586173019,-0.00174278175216347,0.00349570632137253,0.00826738808093386,0.00879950644204519
"2990",0.0104367247377419,0,0.00588883474402446,0.0222890042466346,-0.000438179292557295,0.000695010301897447,-0.00623515977407363,-0.00535924496352547,0.00113396721156644,-0.00186913334812067
"2991",0.00260058326052826,0.00023950493010072,0.000731759623402439,0.00195983038653758,0.0057873935504793,0.00307418122571157,0.0120465293828098,0.0037714014630712,0.00740616905304958,0.0062422403245177
"2992",-0.0169144174466024,-0.00766095219158702,-0.00438755420008141,-0.0134475046697691,0.00278984576515007,0.00148303322623811,0,-0.00214682892751272,0.000432407876689078,0
"2993",-0.018506195510919,-0.0176115548962528,-0.0183621001177368,-0.021561232983661,0.000347678567244269,-0.000197480176524767,-0.0106633146130414,-0.0134480617971161,0,-0.0303970519984572
"2994",0.00340755440184815,0.0135068288006506,0.0153385477487715,0.0184902527711024,-0.000347557728871073,-0.000197214243605082,0.00137868502629024,0.0111778090324917,0.00164262992379394,0.00831735623043794
"2995",-0.00667871690590705,-0.0079960903452243,-0.00368454527516271,-0.0116884161771456,0.00104325125507954,0.000592440599068933,-0.00337919272832965,0.00242644602007713,-0.000776834103427881,-0.0291878088056222
"2996",0.0161443426830865,0.01587691143772,0.0134984481807219,0.012330029070281,-0.00225813418538434,-0.000789683402085295,0.00351619053893049,0.00968265560514392,-0.00112289888026862,0.0045751006142738
"2997",0.00336438248268456,-0.00456834294192809,-0.000912233854500899,0.00695990010606296,0.00113179330239732,0.000987986054997947,0.00312845137563866,-0.000798969282620132,-0.00596681084371165,-0.00390365519694513
"2998",0.0230252252483887,0.0132848760520181,0.0131482406311618,0.0239446858383787,-0.00486928787924523,-0.0000987417246536282,0.00885750513526906,0.013063141209755,0.00374075694843223,-0.00326592898342237
"2999",-0.00218501115761005,-0.00452923865944366,-0.00342450355604973,-0.00867881125388648,0.00393191330440534,0.00256595346393595,0.00136007832557805,-0.0115790613284052,0.00312013355313234,0.00655312555937493
"3000",0.00609537400360649,-0.00574707157870258,0.000904258352552256,-0.000972664391154954,0.00374249757399814,0.00196877888111779,0.00987891704403365,-0.0106497907978395,-0.00172798516896466,-0.00455729637804392
"3001",0.0132414516432389,0.0108381903701067,0.0135525508942627,0.0202044705972819,0.00710028405310292,0.00218598583646723,0.00464654457856239,0.00188391446316039,0.00752988568868029,0.0228908020595362
"3002",-0.0324024227695083,-0.0228735085321919,-0.0369049108196652,-0.0212360533224223,0.0167413748502623,0.00461735034316013,-0.0154575410774033,-0.010475485891893,0.00609912357704245,0.000639377437478439
"3003",-0.00151722494626882,-0.0141429209945474,-0.00148099154787262,-0.00926380561669682,0.00314048451317639,0.00254251560917895,0.025095875955633,0.0114004111835111,0.00017073086994368,-0.00830666140199077
"3004",-0.0232359232203346,-0.00964629347689194,-0.00741563543535884,-0.0187007237741963,0.00186131388579902,0.002926378309555,-0.0141100948009866,-0.00160994713695228,0.00810992836016666,0.0115979115668692
"3005",0.00189718521604942,-0.00774218998111909,-0.00765784318864182,-0.010531709227814,0.00413826774360171,0.000583408072627023,-0.00562689819348139,-0.00833342962212014,-0.00347189443549467,-0.0159236109303792
"3006",0.000226959256249826,0.00352371221984749,-0.000752832345759069,0.00760266234810514,-0.000168240905373707,-0.00252711351632007,0.00073811718191874,0.00135543621911394,-0.00118965839564922,0.00582522978331501
"3007",0.00503556383718751,0.0175569834965958,0.012054954591435,0.0163481719289642,-0.00445825423181823,-0.00272848115506663,-0.0164720117255978,0.0073091418824851,0.00212693549321985,-0.00321752554992527
"3008",-0.000339071844660199,-0.00172537721606758,-0.00297783612273284,-0.000247438493297225,-0.00236587452998627,0.000586214663774065,0.00599927337041173,-0.00322491910039335,-0.00220733506912862,0.0129115793058858
"3009",-0.0184647735061731,-0.0143210179714212,-0.0113870298278249,-0.0141089586810673,0.00347262070073895,0.00156253056480593,-0.00198783224110832,-0.00350500879355298,-0.00399898752658046,-0.0152963551974954
"3010",-0.0196183147934893,-0.00926839021465431,-0.00793042491497664,-0.00928956466038244,0.00582361206836657,0.00292516662311093,-0.0369155092437774,-0.00730518678146697,0.00691957127831144,-0.01165045956663
"3011",-0.00109656381610057,0.000407436689290774,0.00278115888932651,0.00679093340357384,0.0059888366052232,0.00246466855837379,0.00897141187428208,0.00109019812552025,0.00237548988609082,-0.0209561733922374
"3012",-0.0149758370854733,-0.00687370337479176,-0.0147283796344791,-0.0166070966735639,0.0132107576383806,0.00349842405894996,-0.0109535844422687,-0.00490079536413102,-0.00609396519519312,0.00401346090748089
"3013",-0.0162777873691591,-0.00410153153879744,-0.00524157361395283,0.00779414682300961,-0.00363099965285429,-0.00125895060010717,-0.0145928280095525,0.00136813795242463,0.0154134207613046,-0.0093271930529496
"3014",-0.0204895896093551,-0.0123552435510439,-0.0308353699995293,-0.00696042806627306,-0.000165676708239304,0.000872941341168776,-0.0124288750504579,-0.0191255676290493,-0.00436092761423901,-0.00874238444107645
"3015",-0.0264229538174665,-0.0125097244568914,-0.0108739256107269,-0.00934587853935331,0.00497020497787903,0.00251879682820544,-0.0360155714592603,-0.00725838869354234,0.0109501009859325,-0.0110645613123692
"3016",0.0505248578725515,0.0250725692254563,0.0189332452946753,0.0199161497664258,-0.0107154089482168,-0.00473523783137275,0.0327777122568798,0.0187101293747793,-0.00299944183468026,0.0222376880571071
"3017",0.00767746812645287,-0.00411945709985773,0.0133866627396142,-0.00128469012377297,0.000166670594626828,0.00252442217005289,0.00161384634785744,-0.00367326683873248,0.00760484681247364,-0.00951735773123952
"3018",-0.00128999049553091,0.0085315438866238,0.00118288726889437,0.00951889343605172,0.00841387350858325,0.0054238724413127,0.00308806650180826,0.00226885393825937,0.00406401260678435,-0.00823610138714159
"3019",0.00875874190662107,0.00281966718990634,-0.0017723149860307,-0.00458710591541012,0.00379995595987248,0.00375676178115225,0.00307857365409636,0,0.00156948623111663,0.00276814258750346
"3020",0.00104033911451151,-0.00536804788764733,0.00690470967218171,0.00256017091975935,0.00526720398845248,0.0021112656589366,-0.0216171982037157,0,0.000659810309278308,0.00276057124542151
"3021",-0.0238627432606022,-0.00719598153707024,-0.00568181045197358,-0.0181307745701782,0.0113794143746546,0.00794883423600057,0.00641017030720681,0,0.00906616650348369,0.00825877456338286
"3022",0.0334956141325371,0.0300284400703017,0.0338915979776644,0.0322495719599736,-0.0115752152915388,-0.00807607225617257,0.0107060575782811,0.0209396089074474,-0.00808623703340683,0.0136518996195234
"3023",0.00788470144732822,0.00150783918234376,0.00247757272876825,0.00226770469680582,-0.00294814131344379,-0.00277769996239241,0.0100563833234277,0.00277158035790714,0.00345848973223828,0.00740742970686781
"3024",0.00939535904081423,0.00727724970521004,0.0047528428163377,0.00377064596048715,-0.00262831308120715,-0.00249741233623757,0.0181864894889259,0.00801547141772962,-0.00270804199320496,0.0100266691442319
"3025",0.00467353283328498,0.0122074003189594,0.00548729816065374,0.0177811469305245,-0.00156485380703841,0.000577698994649545,-0.00130369024587174,0.00740334007557086,0.00641816017788321,0.0198544006138881
"3026",0.00352746342364596,0.00147669096411773,0.00602180365869343,0.00713586712479963,-0.00643337103178754,-0.000481100059104844,0.0138381382672079,0.00653243194755659,-0.0058866978315214,-0.00259576096476599
"3027",0.000386386731765942,-0.00466944530759072,-0.0115974239925136,-0.0048864049641304,0.00390166266823777,0.00298475551562061,0.0034766039694083,0.00216344479566288,0.00172717334409644,-0.00325304643822777
"3028",-0.00610094564964281,-0.0041974389264956,-0.00359572985025491,-0.00834769879111852,-0.00372102294554566,-0.000575924362045344,-0.0032078641429496,-0.000270114564991486,0.00238089485104531,-0.00848568371229008
"3029",0.0114608710350383,0.00223148755734504,0.0121556742124851,0.00693236750180493,-0.00365215532466223,-0.000960725741985136,0.00991228521495957,0,-0.00172003445720481,0.00790000123072776
"3030",0.00241967099930585,0.000247393852239819,0.00487893649240645,0.0122941095971385,0.000999591388892718,-0.000576810398652206,0.00624611075207149,0.00296908705089205,0.00319986880209711,0.00522536480298497
"3031",0.00758688659107309,0.00519411371772183,-0.00205417860801149,0.00437216802979878,0.000249581984190561,-0.0018277371470975,0.00532046126198527,0.00376736295630864,-0.00130854669113967,0.00064975053065397
"3032",0.0133099310842342,0.0125493199315001,0.0132859960627645,0.00483677285386119,-0.00524144520049485,-0.00318037223025613,0.00378025449498209,0.00294918701151636,-0.00892641054027998,0.0103896539161537
"3033",-0.0135104989292035,-0.0133657815503351,-0.0179132240522069,-0.0173285282966976,0.006774800360138,0.003480507009058,-0.00288716925592802,-0.00534600218597059,0.0035531318018458,-0.00706942989049986
"3034",0.00209248039510324,0.00689662227975751,-0.00282057702270355,0.010286643122537,-0.000415528944941568,-0.000481735327292454,0,0.00618092364023437,-0.00139973655166081,-0.00129445445557619
"3035",0.000531377830543578,0,0.00584572178549769,0.00969699582542582,0.00656582197087774,0.00318113377493123,0.00352506216082604,0.000801324078339549,-0.00156664744035828,0.00259226447945782
"3036",0.00846146006370074,0.0102738747925124,0.0108736453817031,0.0132052185149609,-0.00478908862003491,-0.00230621635189754,0.0116672077933329,0.0122764838675136,0.014617268630515,0.00517138674472584
"3037",-0.00760009264066852,-0.0046004528226361,-0.00723295343790142,-0.0104266858228054,-0.00099553634601679,0.000289018690714515,0.0090525902805807,0.00580022962900162,0.00349991857805709,-0.0135048870193266
"3038",-0.00132709738514425,0.003162290736064,0.000934134022908761,0.00167640775962075,0.00506607043240903,0.00288837469774639,0.00798827351863074,0.0104847252644698,0.00559657713037076,0.00977835680421557
"3039",0.0158308033782144,0.0106692401026993,0.0111981176267182,0.021754736295968,-0.000743688515939422,0.00230422393059748,0.00792486506765511,0.00804169823693401,0.00572672191337187,0.00710137726681648
"3040",0.00878242299186072,-0.00143966380757565,0.00184572243727787,0.00842295418453354,0.0085999436691484,0.00459769627379569,0.0105237975916945,-0.00205875155256152,0.000481177312035008,-0.00512816137458549
"3041",0.000481464905415008,0.00120137918419716,-0.00405301062406771,-0.00788867204345278,-0.00603952458386892,-0.00535084598550795,-0.00682309482801047,-0.00128927826347247,-0.00200400801603207,0.00902057392904099
"3042",0.00703559299879686,0.0028799444735339,0.00221968500880565,0.00163710633152436,-0.0044643033582904,-0.00220931869261476,0.00674932406650819,0.00206557656135997,-0.00433735742971886,0.000638547936024469
"3043",0.00419167662738662,0.00909294683762041,0.00406056674540456,0.0137753520561579,0.0045672663574603,0.00173295980146615,0.00610573001389625,0.00154607429236409,0.00258147791692065,-0.00446711284627554
"3044",-0.00131824599428665,-0.00450556635467447,-0.00827202052250664,-0.0135881702274754,0.000495865542629037,0.000768820590616226,-0.00690153511295599,-0.00617446688455292,-0.00675890736046758,0.00128200777892928
"3045",-0.0095325783692144,-0.0131014247312681,-0.013901771695415,-0.0100396617338997,0.00661004943932575,0.00326525976219405,0.00766829457021889,-0.00310647097681516,0.00243029808116813,-0.00960307277514072
"3046",0.00122142164358396,-0.0036205910115541,-0.00883458626411948,-0.00566050925359562,0.00426822066049226,0.00134013705132174,0.000237961629824257,-0.00103868843867716,0.00379829487309347,0.00129284668618146
"3047",0.000554628732257312,-0.00242247318635835,0.000948170757803402,-0.00332061446599796,-0.0039230614658633,-0.00152963459848154,0.0028529894791669,-0.00285940618554748,-0.00491104584905433,-0.00581019987504727
"3048",0.0128594494930068,0.0109276137047758,0.0176203108923771,0.00832939014270906,-0.00254369858793446,-0.00134032524452898,-0.00580851469767296,-0.000521260066808082,0.00210358417643342,0.00584415558710938
"3049",0.00324673496329697,0,0.00242046825771447,-0.00708050100986224,-0.00378430084385739,-0.00249256386975483,0.00465013762657818,-0.00756398148425075,-0.00395606326533127,0.00581019987504727
"3050",-0.00221810969047254,0.00024020320625362,-0.000742962608969666,0.00190163700867041,0.00569781942297576,0.00470925100941799,0.00320438412100588,-0.00289096861647609,0.00559289116658279,0.0025673722456947
"3051",0.0108972445547948,0.0158500759443467,0.0128252875808565,-0.00142356956944245,0.00156018109283629,-0.000956489437566987,0.00615173150769865,0.00711649524008795,0.00596489611421736,0.0185659623806202
"3052",0.00173064458508909,0.00401902024241663,0.00165172024661309,0.00784030552574144,0.00254114399132477,0.00172350171935842,0.000235021753052234,0.00366392367754842,0.0152243105314669,0.00251418451559937
"3053",0.00201538680668989,0.00565095250040581,0.0010992312621565,0.00565774417866449,-0.00286189074380494,-0.000191116387024515,-0.00705294061777106,-0.00260744006662827,-0.00173633784695348,0.00313475350515446
"3054",-0.00355586992080403,-0.00468270588283959,-0.00146411335623353,-0.00210963338775172,-0.00893876898028223,-0.00296383843668413,0.000828619078213411,-0.000522960855506627,-0.0113061350891966,0.00312495753357278
"3055",0.00619996493848185,0.00305814574866936,0.00219941826476155,0.0110406305881516,0.00595778887380893,0.00297264888771642,0.00532278768389394,0.00313885893985288,0.00359853649903541,0.00249225404025921
"3056",0.00136132425855795,0.00211069496809646,0.00566939857034465,0.0111523657784109,-0.00296131099392349,-0.00152971233803401,-0.00729476816914765,0.00104310828039544,-0.00103583266932272,-0.014916033180699
"3057",-0.000715491178974292,0.00725489906385612,0.00345516241274413,-0.0034466771954148,0.00495005602407739,0.00296816372118403,-0.00272607781640044,0.00442826758244053,0.00167503385957479,0.0044163819462697
"3058",-0.000429444301129123,-0.00348525128702581,-0.00525561257196572,-0.00853122863455436,-0.0113290308974948,-0.00353225181986128,-0.00285242290407872,-0.00440874448217088,-0.00708711566989773,0.00502508265366841
"3059",-0.00186280529286542,0.000932658895962613,-0.00965560334517146,-0.0130232728235646,-0.00340451223903815,-0.00258652324211506,0.00297979102943913,-0.00468876573705412,-0.00561395451737989,-0.00250004222829769
"3060",0.00624387900160994,0.00628940702111547,0.00294329064045051,0.00117813712716908,-0.00924296582763362,-0.00328169588900162,-0.002139069103124,0.00209388915519915,-0.0170175097510687,-0.0112781954887218
"3061",-0.00363735208718352,-0.00416666796219789,-0.00311812862311955,0.00141208152733818,0.00783754239809964,0.00308973119694467,0.00416811302315834,-0.00365638304136973,-0.002625525171288,0.00316865365604024
"3062",-0.0013601674292637,0.002091954792103,0.000919984011975794,0.00987080186106781,0.00209050611093953,0.0005773454451099,0.00308347691750277,0.00550447064830961,0.00131624714241929,0.00505365229360066
"3063",-0.00605690943978621,-0.00185572667612555,-0.00588232820768719,-0.00558539840574235,0.00367149699358449,0.0027898570219147,-0.00484742997249688,-0.00599594230583766,-0.000903713433259012,-0.00565681936947671
"3064",-0.00836550464840824,-0.014640834209391,-0.0118344016466634,-0.0184880609159473,0.00648490265637047,0.00335764929993432,-0.00178234251296294,-0.00131099645446564,-0.000822292567862037,-0.00252848771387459
"3065",-0.00199969133286948,0.000707523013688149,-0.00168415460981863,-0.00715319349546928,0.00421276899850143,0.00143412828397627,0.000952294020167832,0.00709009864997445,0.0109455516262769,-0.000633692099297978
"3066",0.0145011153002079,0.00848454121261688,0.010871684599586,0.0187319824896492,-0.00296124128298458,-0.000763777618581596,0.0147444014764997,0.00547599502541907,-0.00488438635247102,0.00126825226655392
"3067",0.00377083015620228,-0.000934838417954387,0.00241057528928112,0.00518630593197988,0.00701255890870933,0.00277093087266822,0.0041012984045985,0.00233406138060732,0.00605370592365362,0.00633316485474422
"3068",0.00661915296780258,0.0109941885240021,0.00388454321044551,0.00117261114028877,-0.00188420171236703,-0.000381129504531064,0.00455127393395149,0.00569214989053224,0.00699294990259514,0.00629318041424543
"3069",-0.000639710890998124,0.00439610648327671,-0.0106873085292396,-0.00538763571787149,-0.00722324490461468,-0.0014298316671234,0.00151020982473216,0,-0.011547093396224,-0.00437765136383261
"3070",0.00494071857305056,0.0110573163994638,0.0115477232206478,0.0146020521884305,0.00661441807563179,0.0031501065398527,-0.00231982738826642,0.00514531342730828,0.0045747649840775,0
"3071",0.00362566093382011,0.00455690341593651,0.0027619472276974,0.0111419380421767,-0.00057505347560094,-0.00133221016379703,-0.00558088540991664,0.00295662704018262,0.000569244526557489,0.00502508265366841
"3072",0.000248065705367395,0.00362895767333882,0.000367224067863603,0.00045919480299994,-0.00221879278153869,-0.000667027707026313,-0.00292291810563072,0.00179457155750673,0.0027632964664881,0.00250010572949733
"3073",-0.00300990443809879,0.000225887591245533,0.000550624524082055,0.00160630244880355,0.0104603483314418,0.00696026344255585,0.0033421787279051,0.00614099639414212,0.00648405754135339,0.00748116896669782
"3074",0.0112947570299806,-0.00271113613143625,0.00660436383577889,0.00137446093798088,0.0022008985408537,-0.000473306547110086,0.0169491500651402,-0.000762775335334087,-0.00402641327105813,-0.00495051590324702
"3075",-0.0192465171962927,-0.022881754862752,-0.0107526929746663,-0.0292839178927583,0.015534646062126,0.00738917928539795,-0.00601852330921115,-0.0106898281425676,0.00234476875808531,-0.00870642553817436
"3076",-0.00075184613564161,-0.000463794358181224,0.000552653338020903,0.00235682954229377,0.00160180741558125,0.00253904698050156,0.000232851765758602,0.0064316308960688,0.00766312004788983,0.00376411527292286
"3077",0.00745393799219429,0.00417543894801375,0.0110477513066725,0.00305661626897291,-0.00071946657362687,-0.000844282131395757,0.00745054581781801,0.00409013969679917,-0.00496313648676172,0.0018750634218232
"3078",-0.00522903229019478,0.00207900277369832,-0.0034601964802311,-0.0107828494197302,0.00920207480335944,0.00291034531886769,-0.00207999414185167,0.00127289394818586,-0.00522929190918853,-0.00561453565263736
"3079",0.00379060952605492,-0.00437996354663039,0.000548209468230754,0.006635030683249,0.00348862210900203,0.0000936223107586009,0.00868457658811361,0,-0.014152850559598,-0.00313672023395206
"3080",0.00630543831267705,0.00463066352589037,-0.000547909099274824,0.0103577666242571,-0.000948097206681209,-0.00159138250799928,-0.000803622103601631,-0.00127127574897856,0.000902378984374508,0.00062924131247688
"3081",0.0118591626244107,0.0124453407572034,0.012609657522384,0.0165424079595653,-0.0142038715545383,-0.00687625789115642,-0.000344664391682792,0.00305482252042277,-0.00393412828564654,0.00943396226415083
"3082",0.000489727736176393,0.00318692074067584,-0.00685805625158564,-0.00320873483896256,0.00184921293157436,0.00170274995843456,0.00643608041161636,-0.00456841779690997,0.00370282237885977,0.00249225404025921
"3083",0.00157366530471581,0.00816880156406663,0.00599674240995562,0.00689815647109082,-0.0086677104317443,-0.00311628313985357,-0.00102767600928,0.00382452399994948,-0.00147565170989539,0.00124302907589291
"3084",0.0026533352735878,-0.00135055564056674,-0.000541871823048989,0.00616577051179457,0.00283363189132779,0.00104200502215868,-0.00148609649342013,-0.00482597359929382,0.00254513951038238,0.000620774470232011
"3085",0.00484033313966026,0.00157765881058602,0.000722899780049913,0.00771678980591073,0.00129164459527153,0.000473125466911473,0.00686889453381334,-0.00765691331095386,-0.00106459748534438,0.00310163159940502
"3086",0.000762423072869112,0.00180028157779355,-0.00234777321903079,0,-0.00354746531169425,-0.00160788706638071,-0.00591244340512365,0.00282917145326134,0.00434496628107151,0.00371063797274185
"3087",-0.00512498584136034,-0.00539086066455974,-0.00543089582866263,-0.00202705106742251,0.00315552057163182,0.00179988587563318,-0.00480389528771374,-0.00641183600219619,0.00522406325648417,-0.00184842871977575
"3088",0.00341109962147024,0.00338755847421179,0.000181998558285823,0.00473933087900114,0.00241969321111779,0.00236414828558873,0.00907945019307133,0.00877650674160946,0.00308564347404561,0.00864193295515259
"3089",-0.000277505006009759,0.000224972454013761,-0.00309372840647026,-0.0107817377047476,-0.00587384785038203,-0.00226425591023882,-0.00102498392422412,-0.00332664104723235,-0.012790431577677,-0.00489591927758426
"3090",0.00676588510824283,0.00630078789608879,0.00511136584719796,0.00726619820166841,-0.00712248718339481,-0.00463325176248575,0.00524446376355825,-0.000513431956569832,-0.000983968863894291,0.00307492641515528
"3091",-0.00065489367229643,0.000894331420260075,-0.000181601905736906,-0.0051849025071149,0.00252697979586936,0.00133016667173846,-0.00510382407547083,-0.00410987578652333,-0.00188790935093308,-0.0018393001365179
"3092",0.000655322839077099,0.000223498496151997,0.00399637568647071,0.00747787103855768,-0.00626102954395902,-0.00341543748357487,-0.0214317554747951,0.000773596060039461,-0.00896378304216749,-0.00368550360883424
"3093",-0.00244698807359844,0.00402052772631456,0,0.00292402188840568,0.000408950266115982,0.000190474409504038,-0.00908668046321925,-0.00541228784599168,-0.00190858016913809,-0.00369913679082623
"3094",0.00196916897133637,-0.0020022253998031,0.00144742452087487,-0.000672835386063775,0.00523479140072824,0.00237944877129781,0.00681872381479387,0.00155486415716988,0.00074828733578558,0.00309401742611271
"3095",0.000862012736389195,0.000445816278181077,-0.00361334050228201,-0.00650811577890575,-0.00480068555504209,-0.00142431508873986,-0.00980851074627365,-0.00155245030783047,0,0.00493537152270385
"3096",0.00899163110464629,-0.000445617614594718,0.00562100869055659,0.0022588724872199,0.002125801942372,0.00180678326969441,0.0119104780020554,0,-0.00207692941571169,0.00122758060901673
"3097",-0.0022191556279586,-0.00557288773693843,-0.0122611159378654,-0.0135225033359181,0.00815853393703803,0.0037963056992969,0.00652598770128288,0.00207308584016941,0.00291373619096569,-0.00367860027303579
"3098",-0.000616044763689372,-0.00201748556978421,0.00219064128530899,-0.00137088085325665,-0.00145667775530711,-0.00122911680887261,-0.00196826884738066,-0.000775823729397107,0.000830073870423442,-0.00184621621650349
"3099",0.00465672305052611,0.00134763973897556,0.00910750637412527,0.00388933748492981,0.00340385655173248,0.00265067765788052,0.00754055523017971,0.00258809646636937,0.00663517458737672,-0.01171384965108
"3100",0.00156772283371187,0.00471068089012761,0.00397107225475857,0.0020509788130334,-0.00638063200446459,-0.00207725254486979,-0.00955667882626943,-0.00154887197550979,-0.00444921303989754,0.00062387250715612
"3101",0.000510452504931536,0.00468852521263408,-0.00359587334694511,-0.000909732416538689,0.00512116959954301,0.00198713774115422,0.011392694779663,-0.00258530648721444,0.00306211200757911,0.00311710095042761
"3102",-0.00751647175297643,-0.00755557381194549,-0.00342835436595113,-0.00751191561836884,0.0041250329016429,-0.000454448737363555,-0.000689657567646162,-0.00285128520223765,-0.00660061897526276,-0.0031074148247241
"3103",-0.00215899448145618,-0.00425433721474,0.000362104342996439,0.00229358431583759,-0.00476187804341999,-0.00283974540840259,0.000345060810555298,-0.012217153759263,-0.00382059794317935,-0.0112220701642258
"3104",0.00978777893011884,0.00966952893446882,0.0128507441983778,0.0118994028090658,0.00283838110310297,0.00132913138047841,0.00793376813139601,0.0202631696694411,0.0059196263811967,0.000630495656581909
"3105",-0.00411518669084976,-0.00913143646228798,-0.0101858689660194,-0.0205789598319196,0.00274947477448184,0.00255963174296214,-0.00330824592079693,-0.00412706306792565,0.00132611684498762,0.00315068397557128
"3106",-0.0166996765254087,-0.0188806534752602,-0.0182343226885366,-0.0196259817452258,0.00766115219557628,0.00340431491246651,-0.0181984765437271,-0.00207204050787457,0.00331099252232425,-0.0125628342747678
"3107",-0.00138936274545998,0.00504003807611109,-0.00606843938505597,-0.0014130791503687,-0.00432172272725007,-0.00188494071487566,-0.000116507329804505,-0.00285498555870034,-0.00247500208295515,0.00127222146063866
"3108",-0.00302562794052952,-0.00569867301107108,-0.00647540539013314,-0.0158018909141748,0.00409950574697615,0.0026439466827497,0.00233180554777057,-0.00026004311538852,0.00239842023328363,-0.00508254897919436
"3109",0.00502336173633799,0.0066483844030798,0.00689003080324002,0.00599081150444158,-0.00136096904436178,-0.000659284363332513,0.0105850420311515,0.00702933456055765,0.00189771456842536,0.00191564380807363
"3110",-0.0251302789917941,-0.0214074238214267,-0.0225633558986281,-0.0333491113189348,0.00785566557919881,0.00499429208840385,-0.00115104866964322,-0.00646333716263936,0.010211628098493,-0.00509874586703907
"3111",0.00904363778238482,0.00791249180288123,0.0140020005452519,0.014046325565674,-0.00294277516939412,-0.00093758875855332,0.00414845976953937,0.00468384195345228,-0.00171190187840398,0.0134529142144599
"3112",0.00585747899558342,0.00600314713556593,0.00149270465324158,0.00194405215377813,0.00614232254931912,0.00319090795418098,0.00654126244576814,0.000518066985552235,-0.000571615225964495,0.00884951432741188
"3113",0.00926139253582914,0.00895116447166222,0.0040992095080199,-0.00485085013684705,-0.00332990367255159,-0.00196460596533077,0.00592853861705955,0.00569507567809047,-0.00719010545951559,0.00563909774436078
"3114",-0.00646516958760335,-0.00636942136213858,-0.00371129058040376,-0.0180355533973179,0.00222729048520343,0.000468848417466194,-0.00283346833802733,-0.00669244549846948,-0.00707760666484059,-0.00934579439252337
"3115",-0.00661204283768324,-0.00663925184619996,-0.00540138999392958,-0.0042194821409961,-0.00206364309746265,-0.00168660410083987,-0.0147760858910699,0.00492354687087437,-0.0000829092402335752,0.00440255832365777
"3116",0.0090156296829913,0.00691408613603706,0.00692881581097637,0.012711982230929,-0.00159063866456621,-0.00112610512593525,0.00842171704027805,0.00361009021687453,-0.00232093834815106,0.000626152843005601
"3117",-0.00307150571482395,-0.00389105996974504,-0.0081829627278277,-0.00492258566601023,0.00573570476214424,0.00300650442711148,0.00354648399500768,-0.00693722431890043,-0.000997033890021259,-0.0143929485468923
"3118",-0.0122184527851736,-0.0101101873239111,-0.00750040841760746,-0.0128617317508564,0.0112473832493498,0.00608903221479951,0.00136808830168089,-0.000776338753381567,0.00773453106677535,-0.0209523796007606
"3119",0.0022683124419034,0.0106776838857965,0.0154920762800805,0.00100238166212985,0.000861690502552248,-0.000279326591326345,0.00330137242274775,0.00828598784274592,0.00107291410535471,0.0136186761454711
"3120",-0.00930049454034032,-0.010564875485074,-0.0083721113143046,0.00350430742940389,0.00719989981166491,0.00437746242383152,-0.0105525303966989,-0.0118130383131723,-0.00387469899732817,0.00831731624288978
"3121",-0.00671076448656072,-0.009285165666017,-0.00469040353701378,0.00648540514297902,0.00303040284959599,-0.000371000709941449,-0.0119266035558101,-0.000779568854978985,0.000331051885607003,-0.00380710643535986
"3122",0.00273104650859057,0.00585753881111506,0.00452402452182943,0.00545226665115939,0.00859835562829825,0.00361780941748258,0.00406222198885287,-0.0018205939337288,0.00678413981672543,-0.0101910607913405
"3123",-0.0134751884836749,-0.00931751345180587,-0.0106961373725604,0.0034508556212296,0.0125194257448407,0.00665500918533013,0.00416132326378893,0.000260428478920716,0.013476867228583,-0.0263835464521808
"3124",-0.00254292283737911,0.00705399313841748,0.00588009518602739,0.00908876167101114,0.00668911400178018,0.00481150638408234,0.00391396367515329,0.00859607669117235,0.0144328141663372,-0.0033047148998443
"3125",0.0217067013555581,0.0121408250304145,0.0115028899140681,0.00219067259089889,-0.0114014694496759,-0.00366247153001009,-0.0032107074206793,0.00413227943345129,0.000319726638000839,0.00596816962723756
"3126",0.00866230369987786,0,0.000559247266923357,-0.00801550806780282,-0.0056520802949408,0,0.0209363917048839,-0.00411527397145606,0.00255692365070836,-0.0204350464341544
"3127",0.00650248460516623,0.00553645399280267,0.00111802157860419,0.000489777815857018,0.0032261258002082,-0.000183577560316173,0.00146483079235615,0.00335745755006833,0.00326768149145074,0.0174966572558402
"3128",0.0100069309172008,0.0126176168298731,0.0120975126305463,0.0078316013284323,0.00865160934731923,0.00395216629860151,0.00303775027417341,0.00566282545855201,0.00564028453225962,0.00330683328664261
"3129",0.00458905684354716,0.00203887392717506,0.00459726956093376,0.0104420309138338,-0.00941241245232693,-0.00494361894547923,-0.00302855029468529,0.000256025814639349,-0.00995334576043438,-0.00263676074053543
"3130",-0.000242259640459541,0.00520012368932532,0.00329488136825185,0.0112953525142874,0.000613148413860065,0,0.00168759893909853,0.0051176608381609,-0.00119685628027033,0.00660936264706513
"3131",-0.00176530983735024,-0.00584796313740699,-0.0111293988469486,-0.0106939452238819,0.000765640623940245,0.00257591370956578,0.00325733856873622,-0.00865585210275088,0.00519253874420822,-0.0137885081622434
"3132",0.00412623676431312,0.000905040058121198,-0.00110693817028551,-0.00168144473718868,0.00344363430906691,0.00247784720664956,0.00369461168479401,0.00308169280817894,0.0061193355142759,0.0126497765772546
"3133",-0.0011048569846116,-0.00791147278110738,-0.00258585627527896,-0.0110684439992836,0.00251668707269159,0.000732192977052959,0.0016731042742606,-0.00409630957260954,-0.000315955771184151,0.00394477291203388
"3134",0.00038024752332988,-0.000467698857587906,0.00293375329657919,0.00394719683044364,0.00174962175615923,-0.000182877181378327,0.0107165614780229,0.000514091885282841,-0.000632071754615549,-0.00458419598484128
"3135",0.0104709191044263,0.0142722553725101,0.00596243420023201,0.0241758211060821,0.00501149826752378,0.00192142051930455,-0.00177638112897416,0.0066804091635686,0.00506008843152861,0.0118421049993025
"3136",0.00225720160172771,0.00438300432490513,0.00889057583554731,0.00834530156760138,0.00143562539823883,0.00273947288586673,0.00622846648828523,0.00280762079547814,0.00605723711318662,-0.00195051907153276
"3137",0.00955433403224815,0.0101056230765517,0.00973010138533414,0.0146606681790564,0.00264087443286232,0.0016391229658399,0.00442139711163514,0.00763544785308468,0.0251779030821637,0.0201954158937032
"3138",-0.00145348388533384,-0.00159161744179992,-0.00981819195421363,-0.00326268933584439,-0.0109867656013168,-0.00409124461491195,-0.0126554583141408,-0.00303109682148084,0.00663561126812895,0.00255425662399422
"3139",-0.00122454369053182,0.00159415472626723,0,-0.00140287256701155,0.00745654475529389,0.00346904940173043,-0.00624156468944026,-0.000281880681431645,0.0148507808713678,0.00445857696222429
"3140",-0.00980792800311681,-0.00568439378333985,-0.00440685919472805,-0.0103020413273999,0.00309666238281059,0.00154668636303001,-0.0127861348479735,0.00102519334619644,0.00194113032789112,0.00317059845271306
"3141",-0.000997416239863269,0,-0.00147551117842637,0.00946294278569781,-0.00639975876429011,-0.00408787807659061,-0.0188592958492486,-0.00512027237868229,-0.00916539513782555,0.0050568469803165
"3142",0.00354607521523853,0.000228765869366043,0.00406355357645305,0.00703082580433767,0.00704705908941672,0.00300994881146854,0.0115794434933791,-0.00257345191010483,-0.000977701729880986,0
"3143",0.00514568203356758,0.00754453222843843,0.00404710793652341,-0.0013963429297108,-0.000677408835923154,0.000454781315055941,-0.000572445244311659,-0.000257891547153166,0.00271003470972686,-0.0106917812989837
"3144",0.0090786040040356,0.00294984718437985,0.0142909140502754,0.0118852969304599,-0.00233875614736057,-0.00125637813690616,0.00343606244004491,0.00335482750507032,-0.0193693848206319,-0.000635706350688436
"3145",0.00260419536044654,0.00316739058927706,0.00307079620621087,-0.00253331342675633,0.00771335568345788,0.00355549716690073,0.0156375398758897,0.00488679782886159,0.0213597389894249,-0.0165393960464058
"3146",0.00799511469493885,0.00721693661030542,0.00288129605840015,-0.00184724552277449,0.00712898024445163,0.00190756834283623,0.0132613982822281,0.0133094285090061,0.00164905924146463,0.00970239117406657
"3147",-0.00113786963315654,-0.0107478835265966,-0.00430952706425625,-0.00693958302491282,-0.0132628119633508,-0.00634689270613342,-0.0045475578623716,0.00176805208541553,-0.0111502353083054,0.00192190997549258
"3148",-0.00549471074420471,-0.00452691514113779,-0.00577096070937277,-0.00605645743371463,0.00135907261718105,-0.00100364294117838,0.00323135370308081,-0.00353000003284254,-0.00643261697012709,-0.00127885885720846
"3149",0.0012465302129312,-0.00409277634153993,-0.00888806542699261,-0.0030465611281224,-0.000376865304297924,-0.000639504394504886,0.00488669802509079,-0.00328935325050694,0.00350374761616434,0.00320104594039505
"3150",0.00477802070905153,0.00365300231091514,0.00603956233632985,0.00846262446303525,-0.00550691183780505,0.000548427280808284,0.00530489236566734,0.0020309062038506,0.0157874914611007,0.0216975534556096
"3151",0.00234413054232863,-0.00159241021582646,0.00181915544171485,-0.00186482854745662,-0.0133505447481962,-0.00493278838101396,-0.0112136601231343,-0.000253362498208509,-0.00844358501914999,0.000624588412292182
"3152",0.00447704807502047,-0.000455657414430433,0.000363170424888093,0.000700641088742904,0.00115315004333816,0.00110147382612724,-0.00177893730557588,0.000760362643632551,0.00625472508488456,0.00249679418045523
"3153",0.000332632021769363,0.00182362115195867,0.000726058791346462,0.00373386604585724,0.00575932740142293,0.00210930217840555,0,-0.00202598320436076,0,-0.0105851998891362
"3154",-0.00322526863453909,-0.00341302830231749,-0.00743696469138722,-0.00139494950010655,-0.00297731961499192,-0.00219624432208498,-0.00233903118896983,-0.00304481370862986,-0.00846255529440998,-0.0106985729502709
"3155",-0.00680501004557243,-0.00205482098192666,-0.000913770348274223,-0.0030267948703101,0.0107978599463465,0.00467712906418694,-0.00401920310769488,0,0.0164653179667065,-0.00890587338578497
"3156",0.00366089324370855,0.00503319463611973,-0.00256079339209137,0.00607203990052496,0.0000755886346661683,0.00246458847590758,0.000224211230692051,0.00432675665364268,0.014117951937614,-0.00706035519196246
"3157",-0.00555489629853023,-0.00614610619737521,0.00256736789082113,-0.00510682702313581,-0.00234839298110545,-0.00182114300067615,-0.0146812431678838,-0.00405479980500478,-0.0147273963870866,0.00581777724944499
"3158",0.00245643378887284,0.00206134073216435,0.00146338454895445,0.000233249618771136,0.00189831510965366,0.000456130266382804,-0.00181980918838076,-0.0055977828609326,-0.000148761804500963,-0.00321338909511093
"3159",0.00715005715023831,0.00640005437435875,0.00803648435627458,0.00116630967482623,-0.00545694147697873,-0.00164138127258073,0.010141313955137,0.000511531839128221,-0.0056526219186156,0.0064474309978213
"3160",0.00469953596106287,-0.000681415714134492,0.00126829611388213,0.00163101228300588,0.00434348326907563,0.00146145364653205,0.00282010138483058,0.00153469926926109,0.00508634146029863,-0.00448428304224902
"3161",-0.00477717266751798,-0.0104544921902794,-0.010676765512232,-0.00883931988352438,-0.00478008253108919,-0.00173282809499142,-0.00461201136317801,-0.00561801645820514,-0.00707000844943095,-0.00386106898946703
"3162",0.00670002132638436,0.00528251789330536,0.00256084892148234,0.00211223448544939,0.00236366527411525,-0.000182750268347687,0.00339024308360303,0.000513593989693195,0.00164893571651836,0.00129201154218861
"3163",-0.001821190722474,0.00182771844773733,-0.00127714463139084,-0.00187356305370401,0.000304129627502592,0.00091377024515471,0.0029283254876411,-0.00359339600579112,0.00665968277955487,0.00387103320698201
"3164",-0.00245468491153678,-0.0150513285907889,-0.0063938890780636,-0.00774281072390437,0.00243335492774577,0.000456472640067762,0.00718688938309042,-0.00643997968017529,0.00334495654013933,0.00578399589622292
"3165",-0.0109403176062092,-0.00648294383027359,-0.000735421822407156,-0.0122960575234992,0.00804041109103348,0.00255496028101043,-0.00334479196437476,-0.0111486347296466,-0.0131129726807816,-0.00638968965774234
"3166",-0.00870790512363173,-0.00419483324743752,-0.000183953528870129,-0.0196313501550002,0.0198603748446076,0.0113424726365723,-0.00100686143338058,-0.000524480674058192,0.0240221967708476,-0.0276527736668752
"3167",-0.00752960427954996,-0.0100632799074319,-0.00515274518193776,-0.0097680498451983,0.00924141518997446,0.00207362648663412,0.00447931445189709,0.00996862512701746,-0.0038120737830929,0.00132277363287803
"3168",-0.030073047807857,-0.0217492986935625,-0.0247872446882911,-0.0369913456359242,0.01728826131482,0.00863693153997347,-0.0179487374105187,-0.01999995714601,0.0139818530722045,-0.00858656973011873
"3169",0.014022882454499,0.00410817693262899,0.0127085959851618,0.0143406376016595,0.00799316123527816,0.00160564608938385,0.0105573650875894,0.00477067074891946,0.00812839144276589,-0.00532973477973142
"3170",0.000590838815329509,0.00505412797474047,0.00693008501657366,0.00454429455290373,0.0003571969776619,0,0.0104470715392535,0.00501192244569348,0.0151896907295461,-0.0127260991363837
"3171",0.0196199412020854,0.0107759048765264,0.00706851242864848,0.0123146483099983,0.00214241660123737,0.0000890545588685399,0.0167872022537423,0.00524940125948814,0.00503468997206946,0.00542736221015194
"3172",-0.00681151714332895,-0.00497507715621748,-0.0105282273865946,-0.0101788182562097,-0.0019952692673052,-0.00151381970719688,-0.000109392622585358,-0.00365546027843044,-0.0033161716874669,0.00877197552943043
"3173",-0.0121732076425888,-0.00785721171229481,-0.00952025085147989,-0.012039095242882,0.0208496676781165,0.00633184188294744,-0.0038271731313555,-0.00445476794314703,0.00969849956457947,-0.00735781389097367
"3174",0.0155516809162781,0.00863932367315479,0.0113078755944878,0.0126936034863279,-0.00342740283591281,-0.00354477529840425,0.00109761785341145,0.00236906728875685,-0.00595951742412126,0.0235847893992234
"3175",-0.0295676346665993,-0.0271235133822006,-0.0242265731886174,-0.028829206667189,0.0225295511816517,0.00667024496387314,-0.0162280119502798,-0.0168069157522654,0.00684159265652129,-0.0151414293457932
"3176",0.00264177162107604,-0.000244457787457741,0.00954929276952798,0.00671132039367262,0.0111194104022936,0.00636095459251584,0.0110342809693464,0.00988257869385656,0.00665497022767081,-0.00802138964796029
"3177",0.0147549825609603,0.0119862114749407,0.0104048131904593,0.0138462212519352,-0.00801022901580462,-0.00263362379328946,0.00870908978628804,0.0134883867140327,-0.00640221307729039,-0.000673900029193431
"3178",0.0120477980447762,0.0077350491748287,-0.000187191054237923,0.00404646369744643,-0.0143025158644285,-0.00475319721825895,0.00754098704702311,0.00287056979483347,-0.0116963020849999,0.00472013878150723
"3179",-0.00766263661734101,-0.00575667356436949,-0.0020599419144286,0.00201511649957387,0.0103444010561295,0.0044220744469663,-0.00748454618121774,0.00286235321016659,0.00779537943593356,0.00268454096763349
"3180",0.00813555782970377,0.0118213588260563,0.00337778586630177,0.00955249609479702,-0.00666517146263712,-0.00264150826793474,0.00371573694869642,0.00337322072253099,-0.00316441866147987,0.00334674288307091
"3181",-0.000307943346966155,-0.00214587850316972,-0.00149622642837766,-0.0129482152012312,-0.00664080494056507,-0.00220710180899042,0.00555322362031485,-0.00362045631076902,-0.00253951052975143,-0.00466975715446305
"3182",-0.0256872928783553,-0.0126642052673843,-0.0112380586884105,-0.0148839119335499,0.0164345738971272,0.00672435941792338,-0.0137519808200025,-0.00207612413856595,0.0195898452442651,-0.00737260842225429
"3183",0.0110583022777448,0.00701842345292092,0.0145861004558192,0.00537771948421817,-0.00404231731564086,-0.000966745320884588,0.00735616423745444,0.0052014754842431,0.000138752863130476,-0.000675265120282376
"3184",-0.00392362082627495,0.000480624892194026,-0.00317401585972565,0.00178306281537877,0.0154090450063102,0.00431076827816201,-0.00381474864452214,-0.00051753184043879,0.0095707398630871,0.00675673356420781
"3185",0.00704168264847116,-0.000720699816569192,-0.000374598165568285,0.00279675722004358,0.00128716208159907,0.00035037436133134,0.00229757355995241,0.00232981819713451,-0.00281653486490541,0.00872487747592454
"3186",0.0127727989434114,0.0100961790678529,0.00712008917882345,0.011156294873903,-0.00378874203444202,-0.00192644159377409,0.00796852875204657,0.000516624276227562,-0.00716456993208681,0.00266132126566654
"3187",-0.000444126675826273,0.00356969475049329,0.0031627773106373,0.00777320015145233,0.000271436395864688,0.000263264526982887,0.00129965656246989,0.00438807221709103,-0.00256727041934735,-0.0159256794434508
"3188",-0.00584732622070694,-0.00308265942902075,0.000556411697061998,-0.00622041509891968,0.0012925710872993,0.00219643082563259,0.00973384497477547,-0.00565408541858459,0.0139130434782608,-0.0053944247471307
"3189",0.0113505020049014,0.0164129025794546,0.00556070388652974,0.0167751472495858,0.00149438856742523,0.00157798519340546,0.00781915063404348,0.0129232378636057,0.00624359519725548,0.0237287654582146
"3190",0.0128553704353056,0.00514855841283213,0.00718896000714198,0.0113272456274078,-0.0181103080403018,-0.0080524781888337,-0.00627041937292416,0,-0.0240011243965328,-0.00132452568052432
"3191",0.000772105212135443,0.00209551025870502,0.00347728897432753,0.00438284889779061,0.00711514704721772,0.000617558462839618,0.00192505132201659,-0.000765379646751163,-0.00852313125976756,0.00265256475118081
"3192",0.000503457324506185,0.000464656192306956,0.00656573703473406,0.00315151057762009,-0.0177652516448494,-0.00617285049791128,-0.00651155016526628,-0.0022982857597752,-0.00373449131531134,0.00925928103607609
"3193",-0.000234765638702839,0.00139339129405336,0.00289904636497629,0.000724899529996215,-0.0175278563792323,-0.00727585913702933,-0.0106371090616978,-0.00307142153859008,-0.00855793202176902,0.00131050490558815
"3194",0.00711096235810071,0.00533390108254062,0.00885281146502215,0.00700316587316152,-0.00177690447484569,-0.000983311268547782,0.000977458402061648,-0.000256744997346181,0.00606367557744147,-0.00719890871020412
"3195",0.00346370089261216,0.00599775261627977,0.00662602489682618,0.00719429870050825,-0.00655089926242025,-0.0022365808356628,0.00488231900665981,-0.00154078196907936,0.00205635681809802,-0.00395517459858208
"3196",-0.000663749814349246,0.00275165937693567,0.011741671559945,0.00571429432984538,-0.0213590670351422,-0.00914636798876867,-0.0116606258079102,0.00823040809823361,-0.00827917451207039,0
"3197",-0.00308874800530756,-0.0107477833270933,-0.00527511763671229,-0.00781256309453338,0.0127435806797442,0.00434387939318248,0.0102687710597011,-0.0043368013899473,0.0083482914740618,0.0443414722905136
"3198",0.00253191024520727,0.00485441592267422,0.00371219485965035,0,0.00542372936400848,0.00261293333954149,0.0109212425403318,0.00614922249716998,0.00198131181807826,-0.0190114068441065
"3199",0.000598240941616979,-0.000920212368100692,-0.00211345210204517,-0.00405627178753709,0.00424364253876819,0.000359637740673824,-0.0035297153372178,0.000509278051028073,-0.00628530340599009,-0.00645992644230764
"3200",-0.0000664876839169271,0.00345389364657311,0.00741266847814037,-0.00407289001775268,0.00300811986915539,0.000449052219720025,0.00483026970484746,0.00610844683923473,0.00405082774247889,0.00520164843502324
"3201",-0.00472483169611781,-0.00206512466072295,-0.00227751745562499,0.000962295325206863,0.0132107576157718,0.00574723231575347,-0.000427257285982807,-0.000759016138030755,0.0118204842286274,0.0012935513870731
"3202",-0.000234660817604482,-0.00252933908112429,-0.00105352723640928,0.000961345657114476,-0.000211450578842975,0.00142860661126365,0.00149616041573641,0.00104774436532384,0.00559638346826974,0.00258408871869475
"3203",-0.00784682578570628,-0.00576301561431658,0.00140619036464584,-0.0105643026372392,0.0120541768492852,0.00499281458681411,-0.00124670747491573,-0.00357407915147301,0.00528692173913048,-0.0115980023440451
"3204",0.00591477398798235,-0.00486914070573119,0.00403720693090559,-0.000727989074488233,-0.0146270914296547,-0.0065648943369655,0.000753298705972405,0.00358689901245191,-0.0185453815841596,-0.00586701408252943
"3205",-0.00208323769739638,0.0053589206084248,0.00174821624234922,-0.000242864611907589,0.00643251666544908,0.00214323398174487,0.00817204544869221,0.0063824979238889,-0.000282091232008841,0
"3206",-0.00538717378436104,0.000463378343763532,-0.0143105887060947,-0.0128734131819004,0.0024581185890622,0.001425814886028,-0.0060793098356251,-0.0032977380166872,-0.00514842397939885,-0.0039344926789654
"3207",0.00463773963105618,0.00231654147395277,0.00460340617119259,0.00565945449583971,0.00245219735560198,0.00080085313890077,0.00375564550642671,0.00585383953291441,-0.0155253298670827,-0.00987485104181107
"3208",-0.0118947084202438,-0.0108620648461809,-0.00440603555050811,-0.00709559586841457,0.00301044356143776,0.00276940903719836,-0.0105836753385998,-0.00657900464795969,0.00547281650006548,-0.000664871068921102
"3209",-0.017664672843562,-0.0261681867118397,-0.012391625894172,-0.00763931480541102,0.00244326875352985,0.00346324991354696,-0.00388971525908521,-0.00560360530807258,0.0116736370524373,-0.0086494124123877
"3210",0.00819281498589275,0.00695780357436315,0.00501882383157293,0.0129128204795237,0.00912196472917737,0.00522116393332994,0.00976237116141987,0.00768449521225278,0.0045306457783747,-0.00134230457842133
"3211",0.013532119201882,0.00905397540397157,0.0115926782138889,0.00441293463921966,0.00738318913823677,0.00193684962669538,0.00537107195619968,0.0119470162893758,0,0.00806451612903225
"3212",-0.00431472991427562,0.000236196577638292,-0.00634695619869641,-0.00829874887677129,-0.00828825435065661,-0.00333889168665691,-0.00277791175036446,-0.00326543168945359,-0.00852707576576783,-0.0013333559115386
"3213",-0.0155247049744528,-0.0110954095815514,-0.00585524631585277,-0.00713760938652341,0.00269397362218138,0.00211573908669305,-0.00514313183202264,-0.00302422600051233,0.00874259707523506,-0.000667466324014487
"3214",0.00949644004058015,0.00811644237714471,0.00874531607352669,0.00768468867866967,-0.00564865348739563,-0.00255121072227571,0.00323102582478341,0.0050555574234441,0.000916044263191251,0.00267198788324197
"3215",0.00676341876730024,0.00899842411551632,-0.00123852281482706,0.0103320246432104,-0.0148944881744804,-0.0062620369841665,0.00193245076239812,0.00100615527421977,-0.00872935567625432,0.00666220231940717
"3216",0.0103669480498201,0.021121742548367,0.01240040729624,0.0160701558228009,-0.0123768365406983,-0.00683421454620348,-0.000750070102281342,0.0100502236968716,-0.00553937228235746,0.0119126403683329
"3217",-0.00111374381380558,-0.00436681707647868,-0.00437444383659746,-0.00431343189990863,0.00726294222956358,0.00277041034402559,0.000214452551670519,-0.00124378774814637,0.00399912164535543,-0.0045781334059144
"3218",0.00990031926891888,0.0129271410544696,0.0149384778245647,0.00890486456055917,-0.0120883755066904,-0.00481252974225133,0.000536065617439796,0.00697381579263467,-0.00697058843361797,-0.0026280985247561
"3219",-0.00160607914776478,0.000911522426665812,-0.00207797090455231,0.00286263656985342,0.00121642741787875,0.00197007877245747,0.000749982703169616,0.0069255185023307,0.00573026999691795,0.00131747834751383
"3220",0.00294906041527687,0.00478146696455273,-0.00260280208727059,0.00380592940259072,-0.00242979801364107,-0.000357443528350876,0.00556737591749412,0.00147394770685505,0.00142437856493483,0.00394743517647012
"3221",-0.00437713422441988,0.000679757534593373,-0.0019137248191381,-0.00521332050936663,0,0.000894131141481402,0.00798557229001107,-0.000245379913459853,-0.00106673777777744,-0.000655352323614466
"3222",0.0067791575886309,0.00407609380126428,0.00714660775444353,0.0090519864372629,-0.00752259867687077,-0.00366236111463925,0.00728852175246675,0.00588816276290038,-0.00477014072767334,-0.00131149755965509
"3223",-0.00326670353181246,-0.0040595467080915,0.00121149703063694,0.000708128977800593,0.0058471167357621,0.00233100306836942,-0.00325079761788294,-0.000731695515532427,0.00293299964611915,0.00131321984427624
"3224",0.00290951541832518,0.00634054223440583,0.00414868798958046,0.000236028559744694,0.00100462048905081,0.000357659096193341,0.0013675778860851,0.000244077095293393,0.00235379462953911,0.0124589936319914
"3225",0.00163405373209091,0.00360039390117328,0.000516399885898799,0,-0.00200722447926382,-0.000178725048980866,-0.00126077008433645,-0.00390438553301364,0.00711591835989411,0.00518143477574506
"3226",0.00409494961127899,-0.000672616778097268,-0.000516133354693249,0.00707545215445449,-0.00488517308518577,-0.00214627399845146,-0.0102041372330856,-0.00367468916156743,0.00233167527966982,0.00579890297429775
"3227",0.00563650290581896,0.00426287134459868,0.00292641118715453,0.00585476494555115,-0.00909646384594165,-0.00376419371912684,-0.00542021956952676,0.00122951985564179,-0.00860004223459732,-0.00384362468784738
"3228",-0.000296578892536536,-0.00134040244323375,0.00429115214121811,-0.00512228470529752,0.000656060438388284,0.000899681255006612,0.0034195402477315,-0.00122800999297246,-0.00277303045202659,-0.00192926024006812
"3229",0.00306709125989091,0.00626394495282478,0.00273454742982326,0.00444654076114004,0.0146341768219944,0.00485348594791879,0.0055377306062101,0.00442590134208931,0.00549022459893056,-0.00644334190948614
"3230",-0.00266316389767041,-0.00333478382964869,0.000170477625216936,-0.00792161431926885,0.0134901545304225,0.00635060627342066,-0.00169447841647941,0.0034271963400283,0.00999850347472697,-0.0058365754909161
"3231",0.00926384242895217,0.00736111691808872,0.00988411997916749,0.0150304810680795,-0.00307804692209901,-0.00188708512665114,-0.00074266968620984,0.00390332809872884,0.000912764209712646,0.0182648168799422
"3232",0.00401777278081528,0.00465017786621624,0.00674989804278514,0.00994914535714386,-0.0131617353578236,-0.00508341557941472,-0.00775025916468275,-0.00121507343262484,-0.0028760101413583,0.00640612793002915
"3233",-0.00110617942579205,-0.00264493869093796,0.00134096918594984,0.00572734148166232,-0.0112465860933033,-0.00537827115437695,-0.0162636578721959,-0.00364957641106356,-0.0161800077177632,0.00254619201042838
"3234",0.000227969947013351,0.0013259764719431,-0.00217609112971717,-0.00318918141218405,0.00605175887503151,0.00288389941890377,0.00293665847876601,-0.0029303294281704,0.00429024650882015,-0.0107936716004128
"3235",0.00351672874555065,-0.000220766378140391,0.00587145504308784,0.00731274290725459,-0.0181185159663564,-0.00799785141584641,-0.00954335996729794,-0.00269410651361912,-0.0155214884055853,-0.000641891971205011
"3236",0.00246609269730524,0.00022081512669625,-0.000500294710443328,-0.00907444700083282,-0.00420729193705227,-0.0013587525067188,-0.00186133941817068,-0.00982318214053879,-0.00636439556333568,0.00256908653475652
"3237",-0.00190974866623372,-0.00154489809833214,-0.0025029282751281,-0.00709707762687761,0.000667237115588026,0.0010884992435154,0.00230359597533814,-0.00471233197896637,-0.00240192883326229,-0.00640612793002915
"3238",0.00210798550749636,0.00110522832340321,0.00217465200582745,-0.00645605031905561,0.00459251088773893,0.000453086213043852,-0.00700449976333473,-0.00523314937236052,0.00269951120238598,0.000644788954934805
"3239",0.000323653969240834,-0.00198724132789829,-0.00350525584842576,-0.0076584514720679,0.00648881454054173,0.00271714024330727,0.00815608282905433,-0.00551085306508925,0.00400205943399845,0.00193298947981591
"3240",0.00145577214702786,-0.000221214563494887,-0.00435518301594739,0.000701600342905895,0.0103295527507719,0.00505823174645781,0.00798072453541909,0.00428204662978171,0.00420352237146027,-0.00321552085191401
"3241",0.00723638921056291,0.0046470906042555,0.00588838418716042,0.00794580023319202,-0.00108765641414854,-0.000808758682569688,0.00531457542284652,0.00777522534771524,-0.00252591660689849,0.00516131205968251
"3242",0.000737582770329981,0.00132150672653375,0.000836217831834185,-0.00162297612260753,0.00181473693671208,0.00170890225254938,0.00517847885889267,0.00746636159280656,0.00296641327859848,-0.0102695541958202
"3243",-0.000288390845623154,-0.00131976265131262,-0.00317511822330563,0.0020901367221573,0.00833287864266841,0.00188562296589811,0.00128805679299671,0.00370558049468106,0.000505028152684606,-0.00907920528324691
"3244",-0.00371880367307886,-0.00594719046175507,-0.0030175718647133,-0.00440335468351993,0.0103476198377543,0.00367445857690485,-0.000214471015050677,-0.000738385265407038,0.000504672283442753,0.0130890276901821
"3245",-0.00160895214377732,-0.00177270680161112,0.00100883365842619,-0.00209493087638679,-0.00625876841905215,-0.00250023607653149,-0.0137236125641755,-0.00492594986160244,-0.00547704689669382,0.00904394952668475
"3246",0.00222389169582238,0.00244175296572791,0.000671991283627715,0,0.00128810065101548,-0.000179089344335415,-0.00326114352149431,-0.00371291756715653,-0.00188402173913049,-0.000640183169661301
"3247",0.00775018224916391,0.00819308030315824,0.00688260565951326,0.0100303013228731,0.00293083459041443,0.000447690902700915,0.00392627613204133,0.00546591045546463,-0.00479165802266368,0
"3248",0.00226568260957261,0.00109827715633704,-0.00166713796179052,-0.00300232900928166,0.00584421654067446,0.0018794423573012,0.0120587194726023,0.00420046798276341,0.00481472855537302,0.00576553466334007
"3249",0.0044575718486406,0.00153574657871358,0.00200397055985202,0.00115829935875245,-0.00290506935559554,-0.00259037862706779,0.00322018624895337,0.00196863107063683,-0.00529991268694952,-0.00509556275296941
"3250",-0.00370863897235818,-0.00569556505851587,-0.0095000378293375,-0.0157334689917172,-0.00213209634322997,-0.000806141132374871,-0.0027820263153584,-0.00294709195324572,0.00620397073950696,-0.0198463287199427
"3251",-0.00849474360186431,-0.00793127564336493,-0.00201914464399422,-0.000235100245813191,-0.0133329119400732,-0.00359034135652014,-0.0148067971589929,-0.00270928963849992,-0.000507819523372866,-0.00130635779152333
"3252",-0.00670658679760194,-0.00421941390456804,0.00387790695224277,-0.0051727732738055,0.0209674079335203,0.00891816599460848,0.00609880861262813,-0.00197581775610656,0.00957985388677685,0.000654066522213448
"3253",0.00617028885276283,0.00958965082967977,0.0112529604153286,0.0075632594891859,-0.00998516562806484,-0.00383934543119524,0.00389703895082061,0.00222718885591355,-0.00136584716148491,0.0156862734681336
"3254",0.0017979268362156,-0.00176713571407061,-0.00398605851785527,0.00445687497936542,-0.00486409266111931,-0.00233029858802603,0.000862620012036519,0.000987664953866263,0.000575885409960897,0.00193043642338497
"3255",0.00913406893883706,0.00885147598331959,0.0115057535348513,0.00583835770721075,-0.00553457651873435,-0.00305459034545774,0.00172377505000343,0.00666016706235784,-0.00992809352517998,0.00642265108196249
"3256",-0.00314406711882964,-0.004386907386289,-0.00560500436201128,-0.00394700107289137,0.00216822181134724,0.000811023065951488,0.00204340694650029,-0.000980162389044748,-0.00029060457384833,-0.00127634574400448
"3257",-0.00111508034049623,0.00044059931886431,-0.000497375950976875,0.00349648210265263,0.0000722009079927588,-0.00117053145321,-0.00601043923635114,-0.00171697368078882,0.00283470703830924,0.00447288663458867
"3258",0.00283862659765277,0.00484476839009584,0.00215625641740491,0.0146341662473077,0.0078609204243647,0.00414681735399336,-0.00971827344144516,-0.00196562302287173,0.00688553303699702,-0.00445296900902392
"3259",0.00861902015730509,0.00832784148115495,0.0024826298230145,0.0173991890283409,-0.0164579078175378,-0.00790015061746596,-0.0130846452254957,-0.00467752912404051,-0.00352724594770004,0.00894570834782171
"3260",0.00059919623785798,0.0091284730523935,0.00264152806361473,-0.000450028496518762,0.0115676796022472,0.00588180319439058,0.000994318111410264,-0.00296801856868645,0.00447887041358164,0.00506645466891054
"3261",0.00686992229907069,0.0133553244871363,0.00459901053747536,0.00848460659570516,-0.00899017423480797,-0.00467800386022899,0.00642048839211062,0.00620188793447629,-0.0000719884917945723,0.00693133829067927
"3262",0.000219167270232967,-0.00706037624902112,-0.00215626136745295,0.00911985843319996,-0.00137878009011827,0.0000904581587182207,-0.00852816056208616,-0.00665685632262569,-0.000215750873923115,0.0043804543080963
"3263",0.0000625530822258025,-0.00107733247145014,-0.0039893949468085,0.00542254882162441,-0.00821236707915318,-0.00271138271761573,0.0129580399097766,-0.0009927328316508,0.000072002016833439,0.000623031858375089
"3264",0.00409896638667551,0.000215660047117039,-0.00100128508014974,0.000449438202247299,0.0016000209865894,0.000780556667076882,0.00827088089119177,0.00844709515814945,0.00258956257834675,0.00435869731147753
"3265",0.00438418023257925,0.00345050686759762,-0.000668242554823784,0.00202158580413281,0.00131901834100501,0,0.00623426916867253,0.000985475070720554,0.00100444106025099,-0.00123988358548832
"3266",0.00152781651795242,0.0023640662446609,-0.000835840855900938,0.00134492263293162,-0.00146378258838153,-0.000906752090647278,-0.00565216748106545,-0.000157304828414029,0.00308194515246707,0.000252270433905188
"3267",0.0000311515364612713,0,-0.0040154090680945,-0.00223859423499417,0.00285838807968575,0.0017244426733154,0.00273285035744864,0.00262198316102391,0.00943199019861352,0.00441361916771754
"3268",0.00532322091016368,0.00385936972254219,0.00268772052221955,0.00717969486201486,0.0024115661794688,0.00144962936510873,0.00534172763504714,0.00679917009733688,0.00785730139853325,0.00753289391086009
"3269",-0.00024780711309047,0.00384451089278093,-0.00184280452073726,0.00400982410358264,0.0010935945742454,0.00144760363021779,0.00271092123806649,0.00649345456203609,-0.000351193975586694,0.0018692213002629
"3270",-0.00551322197895632,-0.0068085106382979,-0.00889565260504688,-0.00665631240292874,-0.00364109656489708,-0.000632407140381708,0.000756969076948444,-0.00206451431379839,0.00210779874787059,-0.00186573383084565
"3271",0.00242933828322878,0.00599826478149112,0.00321766305195026,0.00223361626088892,-0.00979400102504568,-0.00361597838287098,0.00583535335831864,0.00310328244960933,0.00189293269673496,-0.0062304676779108
"3272",0.00935188367575668,0.00787911004853292,0.0104658841841363,0.0202808116844397,0.0112931826818319,0.00462708504979581,-0.0110657418784316,0.00206230711170763,0.00734781696351927,0.00125391849529799
"3273",-0.00757216073619027,-0.0107754485199473,-0.0110257265114312,-0.0185670384134345,0.0154002062030465,0.0066829323595976,0.00716994310396113,-0.00205806275425324,0.0132685240695074,0.0118973074514714
"3274",0.00381501627650294,0.00363096967108056,0.00354728034548502,-0.00244825283774763,-0.00567845350911844,-0.00107650446523522,0.000862944281291078,0.00232013779146101,0.0104894967058171,0.00185649752475237
"3275",-0.00281180883127474,-0.00574592442026267,0.00168318464904904,-0.000669321731370021,-0.00491579459083291,-0.00143687107763246,-0.0101303823399314,-0.00360080669702267,0.00393515166520908,-0.000617726953815456
"3276",0.0053295821278867,0.00192636982178129,0.000168072598490054,0.00580482237542257,-0.00661093860238493,-0.0023384050667582,0.00239519249330478,-0.00722771690004143,-0.00750152052779929,-0.0148331273176762
"3277",0.0067805937966583,0.00299081386475519,0.00705643481182783,0.00665924543083785,0.00351035611366091,0.000721259733255986,0.000543063188037207,-0.00077999768436543,-0.00565165459858608,-0.00439146800501888
"3278",-0.00287771078399512,-0.00489882843665956,-0.00700699044055697,0.00529221633041765,0.00889087610547246,0.00216186704761334,0.00868428392757803,0.000520386857849164,0.00602619328922938,0
"3279",0.00687735753110474,0.00449484151338098,0.00571238239247296,0.01557356876508,-0.00303387707613423,-0.00116839611263631,0.0106543921821625,0.00546169265449148,-0.00741948791996483,-0.00756143667296783
"3280",-0.00152460103274799,0.000639228638397604,0.000334112924588847,-0.00561550768068053,0.00514418855765597,0.00197965705057968,-0.00383346147196495,-0.000775988593591737,-0.000891544326973026,0.00444444444444447
"3281",0.0022598315594613,-0.000638820286176012,-0.00367403133476907,-0.00781930912642681,0.00663151671537054,0.00251490594432613,0.00887217396420037,0.00336521119599054,0.00583424386252673,-0.0050568900126422
"3282",0.00831838404676954,0.00554014489665455,0.000670482735501299,0.00634853327495621,-0.00315072917329373,-0.00206059636517852,0.00741693961222523,0.00644992298681046,-0.00156950328228833,-0.00127064803049548
"3283",0.00311255687842316,0.00487389287717499,0.000670033489614141,0.00565584064268343,-0.00854817895474858,-0.000807931182548183,0.00115691220103797,0.00410153467573737,0.00184542412474098,0.00318066157760799
"3284",-0.00195815295719093,-0.00801343348854644,-0.0053566118059386,-0.0253082197707116,0.0105056136643549,0.00395326296851173,0.0101901550771279,-0.00663773981492866,0.00109157455189557,-0.00570703868103994
"3285",0.000120729923205554,0.000637733829980336,0.00454394158680382,0.00821125148221813,0.00351341416785456,0.000179007832023848,-0.00571965596806834,0.00411207569417749,0.000340656932647843,-0.0133928571428571
"3286",0.00114685349798638,-0.00403652007648181,0.00117270901612843,-0.0103456086286594,0.00700201846043647,0.00250538270059564,0.0059617114700905,0.00204763080663861,0.00224812327635981,-0.0084033613445379
"3287",-0.0088930892009017,-0.00234643766325848,-0.00384871164152323,-0.0080071398578101,0.00808847341450036,0.00357015813506933,-0.00228743499861095,0.0022988806284967,0.00584557523944995,-0.0149934810951761
"3288",-0.0160293642529677,-0.020525956809921,-0.0179741309923421,-0.0345290822658781,0.0155545275070015,0.0067590566761262,-0.00479359088890197,-0.0127421260311981,0.00682530765847567,-0.0185307743216413
"3289",0.0104791206371506,0.0087316741163137,0.0088949881781557,0.00836035744634556,-0.00783131120464842,-0.00335687473867652,0.00429319569998721,0.00129068699883916,-0.00892678002125047,0.00472016183411994
"3290",-0.000825997901144682,0.00129844192379225,-0.00322141403865717,0.00483655019974893,0.00977924987256662,0.00478646404388217,-0.00312794260478921,0.00567146817642783,0.00541787199193089,-0.00469798657718123
"3291",0.00324535753840283,-0.00129675815863406,-0.00136080963835994,-0.0148980285377487,0.000138381280643696,0.000970331512785583,0.00125506491557958,-0.000256273134421336,0.0000673177928653956,-0.00876601483479433
"3292",-0.0181578801347492,-0.0157974251416886,-0.0163515417535607,-0.020241949744067,0.00912975380378445,0.00502340110191302,-0.0121174520775672,-0.00410258605832581,0.0057924226726449,-0.00816326530612244
"3293",0.00742852226433333,0.000879507475813668,0.00761903030303035,0.0111612678422877,-0.000810041035813391,-0.000851744763572304,0.00306654813657548,-0.00102989114536112,-0.00649568731673889,-0.0185185185185185
"3294",0.0152413054446825,0.0158172671353249,0.0151228907909071,0.0258336765695784,-0.0134670782572184,-0.00580023203782287,0.0102256052068161,0.00489692227095317,-0.0130089511120994,0.00139762403913335
"3295",0.0115480012091473,0.0114618939679112,0.0089723717623158,0.0057234432234432,-0.010934710197444,-0.0043312664690992,0.000208672692488365,0.00051291272677334,0.00122931099231849,0.0153524075366365
"3296",0.0033648125578345,0.00171045542014103,0.00755035260236081,0.000910562258138015,0.00450674377692972,0.000710238232151328,0.0037558725800213,-0.000512649782175578,0.0053883977533018,0.00412371134020617
"3297",-0.00532965351059922,-0.00875131307369525,-0.00965858467374825,-0.0138730949767322,0.0124780923761345,0.00479066773088399,-0.000415780963314294,-0.00461655113184511,0.00264585492452607,-0.00547570157426425
"3298",0.00746532719831561,0.00258402245012967,-0.00117704723092238,0.00553498603470981,0.00276961910400986,0.00194240790734224,0.0100863258690429,0.00566862375160793,0.00257124986804746,-0.00894700619408118
"3299",0.00173306073860502,0.00601372409764345,0.00505048804543806,0.0130733950951099,-0.00504041256158561,-0.00237924760798192,0.00813264128977287,0.00358696812166137,-0.00344195185856722,0.0034722222222221
"3300",0.00644274914880749,0.00576432536293758,-0.00485763810958739,0.0135839263565283,-0.00506594702460472,-0.0025616516772804,0.00796486385129014,0.000510529947559402,-0.000812752246708404,0.013840830449827
"3301",-0.00106696285530883,-0.00785393742615292,-0.00875275206194237,-0.0131784677239224,0.00383625779135266,0.000885518699180299,0.00678748698303822,0.000255302156451975,0.00569345289314205,0.000682593856655256
"3302",0.00160215372147277,0.000855733810195325,-0.00747152330568057,0.000452716161158939,0.00437740020550326,0.00247750703309313,0.00905618861516766,0.00867347377625949,0.00417842687092507,-0.000682128240109159
"3303",-0.00257705863537561,-0.00448907662439235,-0.0148844993176305,-0.00656110844884383,0.00684878491041241,0.00158871157228191,-0.000698014893286691,-0.00354070201387513,0.0128188187919462,0.00750853242320826
"3304",0.00478127256597216,0.00579772385656008,-0.0017367488108111,0.00728763379640163,-0.0000686624354968579,-0.000176291599413791,-0.0125736386957546,-0.00304578472443895,0.00583121712726231,0.00948509485094862
"3305",-0.00410826914499118,-0.00597777540563627,-0.0064370041753653,-0.0156002486999774,0.00783340985452452,0.00290858216604817,0.0108135583992111,-0.0038186503093911,0.00408466320964895,-0.00402684563758393
"3306",-0.0102982407394349,-0.00279211763762632,-0.00840483263167857,-0.00574184644598419,0.00934063281914299,0.00404248879909752,0.00189964789279773,-0.00204456833912281,0.0150252144865768,-0.00404312668463613
"3307",-0.0331653660915764,-0.043291018737885,-0.033727705567231,-0.0374221058576552,0.0149284684553683,0.00778995480061684,-0.0133719272196468,-0.019718350566677,0.00898512622466319,-0.0189445196211095
"3308",-0.0303021989283192,-0.0229625404305511,-0.00164473681204802,-0.00791931883462049,0.00532455968884515,0.00277920719435931,-0.0268028414358152,-0.0107105513683383,-0.0178742588986933,-0.0186206896551724
"3309",-0.00367824356572966,0.000921589819281587,0.00494235758846129,0.00798253507498781,-0.00529635890969682,-0.000519622930146402,-0.0104968109915262,-0.0105623082620163,0.00437050219757662,-0.00983836964160234
"3310",-0.0449116815436744,-0.0303867410310024,-0.0342441153280831,-0.0239980813054035,0.0108486561144376,0.00485270021840045,-0.0524104758003641,-0.0240192858872142,0.000194836655226238,-0.0170333569907736
"3311",-0.00420147991494313,-0.00807217493048862,-0.00113166729536018,-0.00368817328193616,0.0225835950252959,0.011210738124152,-0.031256867405301,-0.0213289247828337,-0.0364934740259739,-0.0173285198555957
"3312",0.0433064746516705,0.0179511732396165,0.0126510954050434,0.0217177196446199,-0.00735747186656133,-0.000683041546917007,0.0481692792348591,0.00558817600221451,0.00552629715843445,0.0227773695811904
"3313",-0.0286324875790996,-0.00893479917551832,-0.012865970298975,-0.00676335716119048,0.0155255232423763,0.0116199851656014,0.000109230753631673,0.0133370250660931,0.0314343303907707,0.00215517241379315
"3314",0.0420330747694149,0.0360615878499839,0.0217227242486349,0.0177528944006053,-0.0106185818058168,-0.00219598975843494,0.0382012643839267,0.0235809889774223,0.00175453246965063,0.000716845878136363
"3315",-0.0332417083933707,-0.0316005739226277,-0.0181179330745056,-0.0210274084123013,0.0248917469047314,0.00888779099776316,-0.021762048698717,-0.00375039898508833,0.0216009400207333,-0.0107449856733525
"3316",-0.0165310908194836,-0.0151335773200856,-0.00960276765952228,-0.0205028064314668,0.0520439069471068,0.0101518520303967,-0.0169800684909724,-0.0188221256761354,0.000380963858627181,-0.0325850832729907
"3317",-0.0780944593433753,-0.087154905778876,-0.0509505722794894,-0.0682781443239934,0.0271031595116979,0.00897010098830942,-0.0741227002826829,-0.0570020271609805,0.00165023798825326,-0.0778443113772455
"3318",0.0517449173722744,0.0360336401893739,0.0298477976701841,0.0508157809792933,-0.0512581064688242,-0.0183569830046986,0.0386113708485316,0.00610284965115615,-0.0211013373183111,0.0316558441558441
"3319",-0.048748479548714,-0.0558517404379727,-0.0338455942423652,-0.0465767868013033,-0.0367976522500375,-0.00997904912744241,-0.0582083324724458,-0.028307356188897,-0.00356035094666884,-0.0180959874114871
"3320",-0.0956771548548002,-0.113471312542923,-0.0980470947472154,-0.100106783238302,0.00619687186364781,0.000508276573690791,-0.0974166748681342,-0.103448218947824,-0.039888262711738,-0.0400641025641025
"3321",0.0854862371124809,0.0606612053181315,0.032812523053851,0.0720854367275419,-0.0226032119315041,-0.00651880893563073,0.085328372185977,-0.0135941605385955,-0.0305162339374359,0.0108514190317195
"3322",-0.109423709430118,-0.113239945289107,-0.0659174194942728,-0.124792477166366,0.0647655626805912,0.0264166645458457,-0.168699975804509,-0.098823558474583,-0.011446119566207,-0.060280759702725
"3323",0.053992088442345,0.0451467268623023,0.0490513408363873,0.0689219749896293,-0.0666830150638034,-0.025072626563892,0.0469908632315217,-0.0193956555662447,0.013555485834196,-0.0158172231985941
"3324",-0.0506329169327246,-0.0688059240975006,-0.0211733348037054,-0.0863650373745922,-0.0564125352426187,-0.013880602504534,-0.0984000761517934,-0.0928109415464308,-0.0199219910827807,-0.0330357142857142
"3325",0.00212493883776443,0.0218687872763419,0.0139702340250061,0.00776950494559747,0.0272255046931094,0.00328149770969888,0.000471100722327034,-0.0612160631446788,-0.0189055014692003,0.0212373037857803
"3326",-0.043094161846041,-0.0126458819714657,0.00244446666666653,0.00738843583001714,0.0751954502261916,0.0254777564612181,-0.043792228132257,0.0236713632580163,0.0149957121484352,-0.0108499095840869
"3327",-0.0255682077067106,-0.00821018035434551,-0.0104190199419414,-0.023915815563909,0.0412093702372403,0.0118347852964105,-0.0505580820623407,0.00334747181113459,0.0441795871516695,0.0118829981718465
"3328",0.0906032620399631,0.0894040036621191,0.0694445132044019,0.0751388083914142,-0.0186144452870993,-0.00680211526389674,0.0800484268339863,0.0930640433246688,0.0485303544388853,0.0216802168021681
"3329",0.0149701792713186,0.0407294808067185,0.0188520519961437,0.0352476450926771,-0.00227125902150904,0.000584640203399545,0.0549027192005767,0.0650602409638554,-0.0136896419956835,0.0167992926613616
"3330",0.058389802701603,0.0487733032258584,0.0328947991960278,0.0378632521279718,0.00492194669735646,0.00242064890990945,0.0741535808558409,0.0282805429864252,0.012822220499229,-0.00347826086956515
"3331",-0.0297856571308275,-0.0345308270676691,-0.00119430727729664,-0.0568439746367654,0.0266927207431096,0.00741118331400026,0.00128363997598568,-0.0352035570223689,-0.00646048660726684,-0.00349040139616064
"3332",0.0324757164586513,0.0187482560570094,0.0121562574730969,0.0164918750519865,-0.00822887264651961,0.00231438982630761,0.0199430350403007,0.00836191593925939,0.00440064367816095,-0.00262697022767067
"3333",-0.0149053853981743,0.000283182332955878,-0.0275645200322007,0.00678463086816339,-0.00811688637184582,0.00181430629333157,-0.0283519281662551,0.00904632457420562,-0.0318466849574507,-0.0122914837576822
"3334",-0.0450048729388943,-0.0467025730708988,-0.0475804423482578,-0.0427777016472985,0.0140105314079517,0.00407130592381622,-0.0659766709788702,-0.0362346283152782,0.00945622405694913,-0.0284444444444445
"3335",0.0230753936154879,0.0190023752969122,0.0127550592526562,0.033670096949501,0.006345863532214,0.000164130342869218,0.00430900257114497,-0.0104650391653116,0.0163934228784226,0.019213174748399
"3336",-0.0144541951756805,-0.0203962995337995,-0.0224600970289693,-0.0189517026946995,0.00237950021251043,0.00073864588820105,-0.015629849352441,-0.0336858976229573,0.00493745904953746,0.0251346499102334
"3337",0.0671662148582439,0.0475907807135867,0.0590508911316299,0.054633200886411,-0.0026112878338278,-0.00451043948646157,0.0750311355862743,0.0381029995946494,0.0277105218883926,0.00525394045534155
"3338",0.00101948204822255,0.00454287323841918,0.0107461070559611,0.00515168875648797,-0.0104724206887115,-0.00444848014209143,0.00970178134091459,0.039437718100831,-0.00535448733571875,0.00696864111498252
"3339",0.0335684148612301,0.014697597097298,-0.0024071816412109,0.0102505982417596,-0.00727604917722091,-0.00124121640448849,0.0715617063719329,0.0202854612965642,-0.00890796630579194,-0.00259515570934266
"3340",0.0152173594687348,0.0239553189997037,0.0130706012467323,-0.00366409244644861,0.00181720883923209,0.00215411770059948,0.0556744639229865,0.0261414212076583,0.0261235574312406,0.0026019080659152
"3341",-0.00913015057670086,-0.0141457026194617,-0.00416838022690791,0.00141454039120448,-0.00912989908174544,-0.00214948745163268,-0.0406947150365636,-0.0071762107220591,0.0171403488923014,0.0173010380622838
"3342",0.029492871225526,0.018763685498693,0.01833769257874,0.0228812698937138,-0.00024413594568784,0.00132563383576545,0.0264305544186747,0.00542103361040835,0.00786809347950945,-0.00850340136054417
"3343",-0.0212481017962827,-0.0392740270462636,-0.00998234488158156,-0.02568351355105,0.0264892401486629,0.00893596716088063,-0.0378523892842125,-0.0287562904385334,-0.00510196112437744,-0.0205831903945112
"3344",0.00482429418115293,0.00281925562956697,-0.00850138361006791,0.00538554437033878,0.0113568978445613,0.00106608166202915,-0.0112405187512169,-0.00740192450037003,-0.000864992244733132,-0.00262697022767067
"3345",0.0270154383300156,0.0334551026145629,0.0133598798261265,0.0222722576184873,-0.0134046566736353,-0.00262144671090347,0.0297739481631336,0.0294556674123789,-0.0194174748876239,0.00438981562774354
"3346",-0.0176179833091343,-0.0136017417628804,-0.0153482683982684,-0.0126861286644308,0.00804484843626518,0.00262833675564678,-0.0362727578537395,-0.0130387898211232,0.00712612694782822,-0.0166083916083916
"3347",-0.0303632484159699,-0.0206839503962466,-0.00939250580750384,-0.0276535761914407,0.0125915639018312,0.0027853198984189,-0.0182736119385349,-0.0264219816513762,-0.00682527251393739,-0.0471111111111111
"3348",0.0221945385300657,0.0152070129657567,0.0173492031470648,0.0272909213648114,-0.0102165921625089,-0.0031043622872523,0.0159744552291834,0.00980022578966366,0.0196708592165005,0.0139925373134326
"3349",-0.0000717269780352581,-0.00776696276746069,0.00138806266111446,-0.00363526306684925,0.00530853507821005,0.000655592892367274,-0.00916048686300919,0.00373266130150562,0.00995486328955342,-0.00275988960441576
"3350",0.0139387063967435,0.012300782778865,0.00772275247524767,-0.00140328371026432,0.00234683170210248,0.000245663743791091,0.00413958873824227,-0.000371885473108402,-0.00428552110409031,-0.0129151291512916
