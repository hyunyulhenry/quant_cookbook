"","SPY","IEV","EWJ","EEM","TLT","IEF","IYR","RWX","GLD","DBC"
"1",0.00212210353361963,-0.0056816367757907,0.010563391559796,-0.0138088934241645,0.00606403628228969,0.00362811560537413,-0.000238385173865874,-0.0074364728506715,-0.01011555892928,-0.0260503050587256
"2",-0.00797640687797585,-0.0147619387360898,-0.0257841292872164,-0.0292383327472667,-0.00435300539131767,-0.00325344210522394,-0.0155036778128443,-0.0124343117072752,-0.0240065523436642,-0.0034512995305368
"3",0.00462554269803039,0.001643580016637,0.00572257607325888,0.00725719426959026,0.00179320457756216,0.000724895474201404,-0.000242365150851409,-0.00338955372229766,0.00515210254785115,0.00519471605092869
"4",-0.000850340852660003,-0.00376400016228162,0.00640098766863351,-0.02233622622841,0,-0.00024134873144499,0.0117533325821724,0.00161926858631745,0.00611769179894184,-0.00861317890472024
"5",0.0033318905730777,-0.00561864703840942,-0.0148410557665737,-0.00230320598256972,-0.00447623771087802,-0.00169152148938678,0.0159282181173488,-0.00565985269618152,-0.00427276924479103,-0.0147698688123383
"6",0.0043803462362455,0.0108136761446265,-0.00502150685504699,0.0126502331889926,-0.00584418263414099,-0.00266348092921154,0.0114344990357789,0.00325279468212258,0.000660191450734482,-0.00132265790941177
"7",0.00759713983333987,0.00905920634572177,0.0129777906266855,0.0203335622338494,-0.00463546913838597,-0.00206333383962631,0.00349645540272192,0.00664595616707353,0.0253999171136414,0.0233996224013486
"8",-0.00195490221031036,0,0.00355838033839606,0.00357474340184827,0.00215913248563493,0.00194650489323811,0.0114984529852964,0.0025765238900326,-0.0032169375331168,-0.0228645994088241
"9",0.000420003593847973,-0.000573262792601392,0,-0.00418511278014622,-0.00306187433362382,-0.00194272337268697,0.00298498396907299,0.00706733772156154,0.0108116506243077,0.00883002834000157
"10",-0.00335620547810744,-0.00305786299936373,-0.000709021861285741,-0.0105519072405733,0.00307127820152053,0.00133798915633787,-0.00343411478717426,-0.00111644408223477,-0.00606642729991103,-0.0105032427762808
"11",0.00196422403411933,0.0107363702976495,0.0070972340763551,0.0179849314068081,-0.00272110489414101,-0.00157883982401452,0.00884496684560454,0.00973966460559961,0.0118856733660673,0.0150376039605462
"12",-0.00308053655416007,-0.00701842472930503,0,-0.00115421535055882,0.00238662142884793,0.00182454767335005,-0.00307384664596078,0.0102783903576438,-0.00444442857142857,0.000871366900456527
"13",0.00294971626693963,0.00897787393321514,0.0056378006431228,0.022753264737692,-0.00657593014833424,-0.00291472791642577,0.00285541522361754,0.00751297955584795,0.0240752866059424,0.0317805604448693
"14",0.00805306403735795,0.00511175045523493,0.0133145224054481,0.0086906108944691,-0.000114456450963196,0.000122564532995861,0.0136674940041031,0.000931827879582681,0.00155688923134556,-0.00843882505047222
"15",-0.0117402398281409,-0.0154452596786125,-0.0165972955541783,-0.0307572256904689,-0.00719064205725684,-0.00389728431586711,0.00595543821868327,-0.00589734210841641,-0.00419717070737846,-0.00893599478055107
"16",-0.000913635159065951,0.00277406200857011,0.000702973492725523,0.00613325054495673,-0.000804167848951431,-0.000121785925859652,0.00301528909831528,-0.00624547015638688,0.00171714023469072,0.0124515654514379
"17",-0.000562763334005512,0.00228931868654758,0.00351369410988456,-0.0132524644959841,-0.00218667529891037,-0.000733636329557696,0.00289490285817817,0.00612762787039611,-0.00623341144564171,-0.020356203459988
"18",0.0052092435246589,0.00532998110438809,0.00630280561297769,0.0154896837802527,0.0011536352728343,0.0009779380324757,0.00344258856019675,0.00405983617508987,0.00705662537243201,0.027705554222162
"19",0.00672329809752248,0.00511180579900117,-0.00417535311128492,0.00775903868721595,0.00840787710839175,0.00366728835409802,0.0113975484885771,0,0.00949861399099006,0.0105308029970261
"20",0.00598248676180879,0.00781804563406929,0.0132771316028601,0.0122480783183911,-0.00120400388486974,-0.000721128708239371,-0.000547244114149303,0.0113528300567416,0.00601571784619104,-0.00375161049023653
"21",0.00138292225767778,-0.000934928409775937,-0.00620668936192759,-0.0030250458743929,0.00126263190095588,0.000856057913550368,0.00711569396240663,0.0110719112766913,-0.0144127872675132,0.0129706315284444
"22",0.000276242655097958,-0.00327417316923606,-0.00763365127702165,0.000953767094085567,0.00137621069935179,0.00110100656062118,-0.000652202644509714,0.00304185694023773,0.000466692602157481,-0.00330437818714768
"23",0.000276239382590582,0.00656985718860481,0.00839182134227956,0.0098735217416559,0.00549673594352118,0.00280726016317656,0.0137045334098473,0.0103103523047769,0.00746389387230284,-0.00497302215289619
"24",0.00220866604647818,0.00372970851324084,-0.000693628373281352,-0.00385933310872055,0.00296201598086143,0.00219291990795756,0.014699868939182,0.00405252116642107,-0.00246957860056218,-0.0120781760068096
"25",-0.00130851508706797,-0.00232218959050201,-0.0124915243617471,-0.00533799804874346,0.000794184139116139,0.000242290864482353,-0.00761365011292536,-0.000598028930855032,0.0137706953630217,0.0231870629732278
"26",-0.00744737633332693,-0.00595934304142332,0.00281112805713257,-0.0119449260115467,-0.00567343629852235,-0.00303652341685323,-0.0141716912726731,0.000598386783463356,0.00915760115190478,0.00618051849681645
"27",-0.0034040630490072,-0.00327846667353826,-0.000700661192873597,-0.00683296171611714,-0.00228186714726553,-0.00133939438962405,-0.0167531470360617,-0.00822136618038116,-0.00680588293379225,-0.0188371198035659
"28",0.00843459960125315,0.00977360148262796,0.0210379789085753,0.0158770136850648,-0.00217363090750444,-0.000732582185716479,0.0178080743151663,0.00813881663311311,0.00258867070469515,0.0183639546801622
"29",0.00656728889566893,0.0128432899816924,0.0164833819574768,0.0215334431225673,0.00951385433666174,0.00573824440902948,-0.00615613543891602,0.0165944620333944,0.00804992454738307,-0.0135245569450847
"30",0.00130471206067106,-0.00202125716209367,0.00810791842247016,0.000594834481790318,0.00295180995688638,0.00157796755879325,0.00825899282312337,0.00294123737616503,0.00060269697441484,0
"31",-0.000479838478015249,-0.000276312491250152,-0.000670054087954175,0.00229403637930714,0.00351081685028398,0.00109069304032294,-0.0034487728589836,-0.00073359923156846,-0.000752943788408844,0.0174491644849777
"32",0.00212713367227191,0.00349948647907183,-0.00335354736799853,0.0026271601940755,0.00225646719954997,0.001210744381684,0.0084360014623841,0.001908258082572,-0.015822829779644,-0.0110249158425911
"33",-0.0004107382914873,-0.00734201954020108,0.000672924936824915,0.00295826191424986,-0.00168897802314882,-0.000121093043859655,-0.00525533507586695,0.0032215221571843,0.0312356463400902,0.0214698305811687
"34",-0.000753266227568772,0.00286605312720845,0.00269009632006356,-0.00252845772484478,-0.00541215398043404,-0.00253984202028479,-0.00506708857912419,0.00627739097785063,-0.00296950268654794,0.013742936552138
"35",-0.00390804618327811,0.00258138706372724,0.00871885215496726,-0.00718182465437867,0.00714264657967156,0.00400094833503295,-0.0141962696164484,0.00681873641717501,0.00848844352975586,0.00637963267720099
"36",-0.000894456295362223,0.00505727465437622,0.00664910159104881,-0.000425567365509361,0.00664051533219867,0.00313999091326211,-0.00648539148583538,-0.00806919656855454,0.00561129643220171,0.00277337747782158
"37",-0.0390578422305794,-0.0539796784832108,-0.0237780825424094,-0.081311219950293,0.0126355050869726,0.00842622641632151,-0.0324191071494272,-0.0368971680434145,-0.0395006472687415,-0.0189648488774585
"38",0.0102508919669144,0.0135397699938606,-0.00135330076077067,0.0250232179307892,-0.0045278005210635,-0.00346168899587496,0.00777621075722745,-0.00558101754437623,0.0163583387030521,0.0153039919303792
"39",-0.00298006655709948,-0.013167931062622,-0.00474245081244884,-0.0143761564979578,-0.000633749723080279,0.00090178533373253,-0.00624079652560627,-0.012133598345716,-0.00992784251228152,-0.00713994426755238
"40",-0.013095321162951,-0.0130538961058958,-0.0163376808281281,-0.00926532892369736,0.005013388265942,0.00324212490240439,-0.0206669344545281,-0.018885825341054,-0.0320571406867212,-0.00918906513063011
"41",-0.00951861568431156,-0.0202800765651187,-0.014532936583849,-0.0256479622984717,0.00166296163279633,0.000598757833027985,-0.0354437051069167,-0.0228478056614959,-0.0122429604809757,-0.0149191936410714
"42",0.0171088805730706,0.0276002293848976,0.0238764454133826,0.0439037548308574,-0.00298843876183408,-0.00131612673416148,0.0344498595743716,0.0281869730822666,0.0193866518353727,0.00941465989397505
"43",-0.00100171391974091,0.00194610296908548,-0.00205764946924714,-0.00609930569135919,0.00388528945902333,0.00179653989211603,-0.0142558194398474,0.0118380434471714,0.00233828519600054,0.0137874316339257
"44",0.00845540241252229,0.0103924539652287,0.00893483065341782,0.0258289395898543,-0.000884456791262478,-0.000120041862419984,0.0160030866019889,0.00369442672213816,0.00279937778540984,0.00160000109706515
"45",0.000284015066560173,0.00288361878646293,0.000681175979498017,0.00178600345301949,-0.0105141116898361,-0.00561925403503527,0.0122499036556738,0.0111961544792041,-0.00356704387870443,-0.0131789655455684
"46",0.00149125909727643,0.00383421155197872,0.00816888225384349,0.00490170329167516,0.00391497552660192,0.00276474062086041,0.00507178047660184,0.00712903990622649,0.00186775097276271,-0.00930789262729326
"47",-0.0194335762900368,-0.0244438542772334,-0.0182309954562265,-0.0290907922056569,0.00601625551626084,0.00443734566893839,-0.0263757925991136,-0.0191262861944046,-0.0100979022791097,-0.00776139923920816
"48",0.00745042423621611,0.00371948082382878,-0.00894089033786849,0.00822154107319983,-0.00454093876928752,-0.00131297752199422,0.00471110692093468,-0.0196534118862111,0.00345257370601737,0.00205841743606472
"49",0.00136349562667348,0.00477789285712404,0.000694109827551914,0.00815421392126936,-0.000111362488093625,-0.00107580534318608,0.00750261759556059,0.0117463042588273,0.000625602136778314,-0.00616274323701982
"50",-0.00279950923513195,0.00349382276014798,-0.000693628373281352,-0.00853779652473619,-0.000222293327685419,-0.000119586210901024,-0.00558485362655015,-0.00346399559345412,0.0100031728665209,0.00248040983341546
"51",0.0120551426129676,0.0149903932102602,0.0111034753177173,0.021936340560097,-0.00211549431888813,-0.00131723366529901,0.0100630547806304,0.0194856548840034,0.001856932751922,0.00494845688755019
"52",0.0054916707618804,0.0098141898189017,0.00892233284910593,0.00656379854202838,0.000558314659723225,0.00143872932146971,0.00324407499408674,0.0151371857308402,0.00818657733044725,0.00123089067396864
"53",0.0164578084874962,0.0245330219404345,0.0108843439286357,0.0299608459278142,0.000446412656245121,0.00143577292448027,0.0140869873044263,0.0227445661451007,0.00842658227791837,0.00163947728165459
"54",-0.000767959612961278,-0.00653898905329087,0.00134601531817791,-0.00427774520985602,-0.00791156661671233,-0.00334572469525696,-0.000796544058840776,-0.00589086577830722,-0.000911546642357819,0.0163664913648924
"55",0.00146678836054392,0.00519143427829727,0.00134397881587867,0.0046398869887041,-0.00280759748095671,-0.00155930137164839,-0.000264295727833486,-0.000444485447961607,-0.00927615543564009,0.000402619932218462
"56",-0.00132493054749194,0.000737474612676925,-0.00536931859607703,-0.000598548431897439,0.00123905029449745,0.000840777048616959,-0.0155083867379672,-0.00340888750680213,0.0105908515551543,0.00442656260043939
"57",-0.00237442375332653,-0.00608229198296961,-0.00404840644282045,-0.00445031885248581,-0.001687279188479,-0.000239854354311397,-0.00828464388015993,-0.00654346572507636,-0.00212635189102994,0.0028045321486756
"58",-0.00727982618867917,-0.00917947793495455,-0.00745257439878999,-0.0178803108458166,-0.00202828377450004,-0.000119930704086335,-0.0116483998518214,-0.00748472984536486,0.00532733662073093,0.00958850037405323
"59",0.00105750355603229,0.0103874221172522,0.00136507899082283,0.0198688581471615,-0.00135460573927904,-0.00144085595347188,0.0053573062485841,0.00829491269040239,-0.00605603303303415,0.0193905524746216
"60",0.000211525865879914,0.00342677556692084,-0.00681640467845968,-0.000171355396247574,-0.00192279016419283,-0.00120192329978308,0.00935415206862622,0.0127148980181369,0.00137084535046927,-0.0147516879941152
"61",0.00112663199934038,0.00360023962951761,-0.00549084484103757,0.00686664768907619,0.00166001141863426,0.00111194907220247,0.0118495498510547,0.00531777099806963,0.00167325834113963,-0.00985019969883938
"62",0.0107629421344138,0.0129677674468172,0.0082816349732866,0.0163682805035688,-0.00124800956511806,-0.000844545217002834,0.00869560182261786,0.00573038101891399,-0.000303659842176507,-0.00397922538928086
"63",0.00111331672350024,0.00254205554440734,0.00752923624342805,0.00629075731786122,0.00102198837922818,0.00157003439987458,-0.00655194861057173,-0.000876957972832493,0.0148867684980474,0.0111865837697289
"64",0.00271116023534979,0.00443765746700975,-0.00271748746451528,0.000917168939095214,-0.00374579073080195,-0.00253362154467429,0.000809585479322861,0.00438692379958261,0.000748435885299825,0.00197546276217331
"65",0.0013865610845718,-0.000991783741184027,-0.00136254036625527,0.00574628847387038,-0.00661030020430986,-0.00459370984506446,-0.000693636421391197,0.000145526353868997,-0.00493571634855339,-0.0102523310478511
"66",0.0011768146455029,0.00722039235042771,0.00341090420667567,0.00471949025603746,0.00298407181082228,0.00206513221264215,0.00254516532846094,0.00611395457059905,0.00946948759160504,0.0139442326305543
"67",-0.00408013520420347,-0.00394268702466438,-0.0040790961759759,-0.00923019103917688,-0.000686924082561768,-0.00121276417532412,-0.0133854380699031,-0.0111404952092401,-0.00119121493798613,-0.00157179448515576
"68",0.00444389738531714,0.00710679998609454,-0.00136491117473481,0.016719533524002,0.000228467956290723,0.000971348721768628,-0.00526295594420523,0.00555969941190781,-0.00134174116452757,0.00590315003881492
"69",0.00456243731490313,0.00741407490509571,-0.00820246670982772,0.00490876933634854,-0.00308923365980673,-0.00169682199447663,0.0109351229707519,-0.00334627609187088,0.0126884314879365,0.00547739648670853
"70",0.00949589765799952,0.0117040134478787,0.0144728618643819,0.0118862491695757,0.00550895668721529,0.00109321469619017,-0.000233184478766857,0.0157660463727354,0.00825480591125038,-0.00778202330855171
"71",0.00265890408237723,0.00131487741645953,-0.0061140701715745,-0.0053909414240072,0.00559411679272692,0.00424531125120087,0.0143095109809188,-0.00546109897937164,-0.00584798228514671,-0.0101961268708496
"72",0.00122397487806736,-0.000525239272527012,0.0013667767035308,-0.0074419580285866,0.00499500875446235,0.00229522301857932,-0.00355612204971456,-0.00173405956055872,0.00558819117647058,0.000396154335922549
"73",-0.000272057327716957,0,-0.00477812258856147,-0.00806817275246119,-0.00169474262004798,-0.000120020401279564,-0.00863241204372656,-0.00376390423506989,-0.0124305065412623,-0.00277227922738532
"74",0.00944108720459624,0.00796914864706655,0.00411529893849427,0.011913168259081,-0.0026021615731141,-0.00108472470608645,0.0109139565326841,0.00624842802153558,0.0173256036920717,0.0138999306258629
"75",-0.00376799533801808,-0.00564721918922007,-0.0109288878774797,-0.00397848233731102,0.00363052654947271,0.00205064557544876,0.00849893308917271,-0.00216629379295341,-0.00640458543251454,0.00665883749617335
"76",0.000405366198928503,0.000174677547557733,-0.00138150846232821,-0.000162956626650002,0.00372939442339448,0.00192678211154784,-0.00683333088181226,-0.00723592452552824,-0.0077644152427655,-0.0136186866940441
"77",0.00918155172750246,0.0105702804708618,0.00553270105156156,0.0123928047805584,-0.00349093628557173,-0.000601062221885273,0.00137619569478686,0.00918416853502046,0.00236226181770594,0.019723922310988
"78",0.00113760350112835,-0.0031116742425229,-0.00481435483137005,-0.00265767907664238,-0.00723211291253301,-0.00288599723782879,0.00137377194383959,-0.00548934738281359,-0.0150242453236743,-0.00696329557888986
"79",-0.000802250316934705,0.000259844150835908,-0.00552855810387898,-0.00500643448901328,-0.000227099078244919,0,-0.00331553868336554,-0.000726146419039786,0.0103184532532472,0.00506419748851039
"80",-0.00829247792945154,-0.00390097414159474,-0.00764451636393459,-0.019314716257139,0.0104741963136343,0.00434150021576007,-0.0191601799755469,-0.002180139824003,-0.00695680896852591,-0.00891469419041446
"81",0.00256263859902117,0.000260977068434975,0,0.00397194030411385,0.000723440941364117,0.0000489490711585994,-0.00526403279765497,-0.00335029292605882,-0.0059620513317663,0.00195550177609105
"82",0.00585213318737865,0.00539455913664466,0.00560244127244647,0.0198646659735173,-0.000565060868801925,-0.00120617154840141,0.00823122054606285,0.0201694784778645,-0.000449812552112516,-0.00780644828912236
"83",0.00541666921303174,-0.000865359537565835,0.00139281789790369,0.00840559396352991,-0.00226097567143868,-0.00108576867143484,0.00396543312744924,0.00286537159367262,0.0124511543683676,0.00472082218868608
"84",0.00379092108247714,0.012126463475308,0.00347729780502304,-0.000320648101281185,0.00407957347480425,0.00253735162495072,-0.00499524159339337,0.00628566769156058,0.0103719665245805,-0.00195784038455937
"85",0.000198711242331617,0,0.00485049973413054,0.0064943803734796,0.00270915909848446,0.000844001015591678,0.00093383894627963,0.0052528563014298,0.000879865057050289,-0.00470760579377849
"86",-0.0013248651740253,-0.0089859063691422,-0.00206876928986777,-0.0129839880546897,-0.00225155828598878,0,-0.0065320796537951,-0.0121453051920888,-0.00542128937728936,-0.00630683405612698
"87",0.00271948452287707,0.00276368589957077,0.0124394946607145,0.0161403792744812,-0.00394893576359823,-0.00325236406853091,0.0116241067748695,0.00114352895486602,-0.00633470858874685,-0.00515664530307158
"88",-0.0104521844666897,-0.0201518346802669,-0.0150167289565023,-0.0244615604206458,0.00237942121197832,0.00253770247141016,-0.00998138420626915,-0.00756828701949352,-0.0214973619643007,-0.00398732915969924
"89",0.00855709188815768,0.0168744201175179,0.0076227493308112,0.0254005169329854,-0.00350316973415132,-0.00204836075805004,0.0111372896401729,0.0141007231080379,0.00681813636363637,0.0148119473263204
"90",-0.00218726938167213,-0.00216051656050609,-0.00275127729948732,-0.00992443693385447,-0.00260732750316151,-0.00144907312466036,-0.010435057630942,-0.00397277154726183,-0.00255828453987728,-0.00355029840873888
"91",0.000265430626462004,0.00259840518395249,-0.00827560700992136,0.001203018863837,-0.000341363628788227,-0.000120547120370129,-0.0134741148694317,0.00284916056142892,0.00392278219557607,0.00989703519012286
"92",0.00684100533329213,0.00216025800250552,0.00208618207096434,0.0144975677307329,-0.00068270311463936,-0.000605315762566061,-0.00926381233148488,-0.00724444091890808,-0.0141268858712521,-0.00980004381165411
"93",-0.00197917191097019,-0.0017244707161066,-0.00832761181988406,-0.00363204127471539,-0.00409687162839201,-0.00266206243198097,-0.017981289059617,-0.00887118914632656,-0.00823170756803993,0.00831350277362031
"94",0.00872502712514911,0.0125216096633798,-0.00279908790985928,0.00515061126853289,-0.00662784140795758,-0.00291204364921682,-0.00866652095420395,-0.00389730532460486,0.00707038140394678,-0.00157051832110122
"95",-0.000524842444591611,-0.00759063781014657,0,0.00181359499783329,0.00299038865978862,0.00133945534178292,0.0068954709459379,-0.00130481947198891,0.00228939265671824,0.00983104263365253
"96",-0.000786334689572454,0.00120321445642357,0.00982466261917581,0.000157116156886294,-0.00516128672913585,-0.00279510510024372,0.0103953583586696,0.000580921952685332,-0.00715701255236845,-0.014408109306017
"97",0.0001315707318994,0.00472094955185298,0.00138974315944718,-0.00157363334664318,-0.00288174957659115,-0.00195046014050526,-0.00786769094037953,0.00203027227571084,0.00521478551601784,0.00474108523167938
"98",-0.00905329253452414,-0.0105936811341796,-0.00485763849449883,-0.0240349429496579,0.000925432505557433,0.00134311695463429,-0.0152494408648298,-0.0123029817097307,-0.0120537227333885,-0.00550522883832627
"99",0.00417075139750245,0.00682163001474634,-0.0041844095016087,0.0153415333315705,-0.00231101535320954,-0.00109708971648625,0.00631804507859823,0.00029329796809896,0.00293439382239402,0.0122577335130811
"100",0.00362536810744873,0.000428654478512813,0.0105047118891903,-0.00341967397596821,-0.000114829211280032,-0.0020755568959433,0.0305307325965118,-0.000586098115259337,0.00200181700025182,-0.0218748918446232
"101",0.00814506343286747,0.0048864426121269,0.00207854829292375,0.0102137958040429,0.00208384116807303,0.00097902247651005,0.0255641737553167,0.00630326419324367,-0.00537880743814345,0.00958467109811956
"102",-0.00104184770089621,0.00153558899638284,0.00968206744539613,0.00284365313684387,-0.00184874958620462,-0.000366778599781403,-0.00267890408319782,0.018062406561407,0.012669962721416,0.00909802267606286
"103",0.00495673347246339,0.00894352709682789,0.00547949940028669,0.0249687210202629,-0.00525359330742337,-0.00430833778719675,-0.000467042864799927,0.00300471002029967,0.0137320870654245,0.00744810721222477
"104",0.000129563533615373,0.00303969311022922,0.00340592176576959,-0.00445693920652723,0.00455680856270058,0.00160301607518099,0.00630969501976941,0.00699056402063847,0.00150510230267598,0.00894950605841682
"105",-0.00395841371612271,-0.00547105332597608,-0.00135758160328481,-0.00347400234196626,-0.00628095196194711,-0.00320023578512063,-0.0173013004456121,-0.00878355773901729,-0.00255482412752006,-0.00385662185426483
"106",-0.0107501220507022,-0.01980371933167,-0.0040790961759759,-0.0251740433300561,-0.000467774431446744,0.00049345206141882,-0.00626243788333136,-0.0195799319777034,0.00060269697441484,-0.00038718847866448
"107",-0.0180453456611517,-0.0231393388972323,-0.00409538381154551,-0.0154151495817942,-0.0179155396202174,-0.00999608375027294,-0.0309158365935657,-0.0236151323284872,-0.0173166982492577,0.00503486046064849
"108",0.0130118891383362,0.0142301856684051,0.00479760279730379,0.0176741313747513,-0.00083469885408749,0.00186974068483181,0.0164413734427369,0.00104487271594467,-0.0159362698150086,-0.0177263688049796
"109",0.00172104257570549,0.000435722407928774,-0.00136412690040255,0.00856431627366128,-0.00286352649258126,-0.00261295873015166,-0.0147264880476032,-0.00372796120775742,0.00747424466717161,0.0192232805596453
"110",-0.0109052656036537,-0.016463364007074,-0.0129781881742825,-0.0173768535828651,-0.0144812901542792,-0.00711026470811182,-0.0210732940271374,-0.0176644394547724,-0.00927355529861917,-0.00269446454548161
"111",0.0149682234660333,0.017270416078762,0.00276811560760759,0.0200051817306981,0.0119000405423866,0.00326630393594796,0.0215269375108065,0.0118865398930532,0.00670828414066427,0.0127363633446651
"112",0.0063862773713439,0.00948969811085609,0.00138038560829989,0.015689359443515,-0.00251980271872465,0.000250361378528963,-0.0102915758348973,0.00135499807753425,0.00108475129528518,0.00952748724430674
"113",0.00568988631004275,0.0125054105713351,0.00895931201158828,0.0227856209871451,0.00685751157967895,0.00438230983648946,0.0151026194995756,0.00811284466027429,0.00386996916006099,0.00604001949708444
"114",-0.00117615517240899,0.00212933320753894,-0.00204921633145361,0.000905838168359541,-0.00203126353301342,-0.000498257730639939,-0.0148779238763278,-0.00330946061417603,0.00154200467361609,0
"115",0.00248559790887759,0.00144523061509472,-0.000684460724354352,0.00113212468296653,0.00933935031738886,0.00486362818036623,0.000990073237193245,0.00739523711683621,0.00816021592733862,-0.00975602421892541
"116",-0.0138975330591123,-0.0129860345427952,-0.0068495479033589,-0.00851659163164475,-0.00806632952175035,-0.00322673092937631,-0.0178083981384648,-0.0112362440008836,-0.011759376370218,0.00113671378480618
"117",0.0055575929902314,0.00610535300503789,0.00482787013365482,0.0124663313011013,-0.00478347008885871,-0.00124543027134205,-0.00402977970359808,0.0037880988384007,-0.00231804979629191,-0.00454197639049791
"118",-0.00940881712618946,-0.00965815088848165,-0.0096085671741567,-0.0132133396071092,0.00648904275201589,0.0029921136764397,-0.00379242182721107,-0.00981144665042721,0.00340769837074673,-0.00228145187285711
"119",-0.00478195195278541,-0.0027617052255775,-0.00554411585060943,-0.00760807049348711,0.00549188947205215,0.00323145784554169,-0.0227155119529341,-0.0213410321894127,-0.00540288677682743,-0.0038110602241177
"120",-0.0102785739490165,-0.00519239127503512,0.00139361690690842,-0.00873986715170738,0.00023638320707442,0.000248071546815387,-0.00142854615881738,0.00233659557967791,-0.0125717988514669,-0.0114765510385546
"121",0.0142289351664922,0.00913461583706021,0.00208763378414978,0.0142308411082699,0.000950160039906667,-0.000123644481701546,0.0217164748829937,0.00310765801925594,0.000785900672522821,-0.00154803023238326
"122",-0.000132826643915895,0.00206876905301168,-0.00208328464873508,0.000228542657458419,-0.000236993827898324,-0.000619689643849508,-0.00390631293038701,0.00898523256849959,0.00926659366315663,-0.00310073611494466
"123",0.000332075846521063,0.00593619782948629,0.00974253336449094,0.00350692260469398,0.0103194807524911,0.0052066724287787,-0.00128975372707874,-0.00230310842972414,0.000155539988934361,-0.00077756390523942
"124",0.00904066314606111,0.0116307451768884,0.0179184334085294,0.0202841510689635,0.00525685190679592,0.0015229525480227,0.0251872710070575,0.011080236238143,0.011669519760519,0.00622568534584866
"125",0.0036235085168721,0.00608661609766581,-0.00203101387778337,0.00796746331164333,-0.00609648593953283,-0.00296756591706804,-0.00466145689999586,0.000456887969964903,-0.0043063520904193,0.00116001076655725
"126",-0.00105025194418706,-0.00344523687316478,-0.00271371736058579,0.00443223016955163,-0.0112070217429092,-0.00557821620424104,0.0160755470365697,-0.00654184200317254,-0.00494284846904058,0.00926999570093279
"127",0.0052568668248314,0.00758873382578495,-0.00476164045462701,0.0171358553490217,-0.00405577024203163,-0.00236884264990844,-0.00211765383904794,0.0124041656952312,0.00838250569334065,0.00841948881502264
"128",0.000784367934051344,0.00343090861921747,0,0.00968932290718083,0.00359303157530588,0.00362407264998565,0.00374535631760686,-0.00862187604070552,0.00646548655273227,-0.0022770415146578
"129",-0.0142386324486269,-0.0146774293747713,0.00205028058654677,-0.019693618826147,0.0169497447334273,0.00684773618236245,-0.0304727500752756,-0.0122063099249407,0.00351795672306299,0.00722704709078603
"130",0.00708968087496209,0.0131184605122894,-0.00341054784073358,0.00825474566485651,-0.010329123239225,-0.00346216034776159,0,0.00447930672792429,-0.00259105315361896,0.00226594368689348
"131",0.0157905196546597,0.0167085826590549,0.00684479655351522,0.0219534080641952,-0.00343822002851113,-0.00285419058380276,0.0125721485655106,0.00830393358407311,0.00886300400785434,0.0026375300692274
"132",0.00297901582226356,-0.00246503612406057,0.00475854860120717,0.0124068966361972,0.00273686714722388,0.0022403814940839,0.00950176623026699,0.00732044809283461,0.000151499552476508,0.00150315505542631
"133",-0.000129136619286707,-0.00230627679613626,-0.00202988876365118,-0.00980407953931961,0.00961316143634194,0.00397260276321121,-0.00552180265466806,-0.0040880759013282,-0.0031803574614625,-0.017636035275769
"134",-0.000516096611510641,-0.0013211846764013,-0.00542383856701623,-0.000777638964366001,-0.00211642564650216,-0.0021025704374843,-0.00643603504540946,-0.00881734388375843,-0.00106350653296861,-0.00611145817995895
"135",-0.0018096814027867,-0.00727512271277853,-0.00477146232650705,-0.0122442839600722,0.00376940582558638,0.00359509632742028,-0.00546131296624808,-0.00153344991013771,0.0132319847908744,0.011529517868204
"136",0.00388431530809896,0.00441373909893872,0.00479433833123522,0.00995977460861242,-0.000234217999210751,-0.000123194316603681,0.00331976069663442,0.0015358049901617,0.00585408259438247,0.00341949609782533
"137",-0.0101245258600619,-0.00920313982412357,-0.00408980091024624,-0.00688172231123785,0.00903838997340212,0.0049406410758015,-0.0160378540429779,0.0007670632748773,0.00850619285162812,-0.000378725846339356
"138",0.0030617879056456,0.00317977636782385,0.00616010445030502,0.0289328116681262,-0.00162863299338367,-0.000368778517039314,-0.0174648254695839,-0.00766254063832905,-0.00162771525221317,-0.00454541746867632
"139",-0.0173411411754499,-0.0212710353126748,-0.00340137185034006,-0.0342293707330035,0.00372881926361601,0.00270515279194594,-0.025674854722873,-0.0200774394506253,0,-0.00761027412690252
"140",0.00204922760069404,-0.00196080239206564,0.000682570960927942,0.0057514560287284,0.00197323246120029,0.00134873264824686,0.00135119606680845,0.00315237138009361,-0.00844818425302818,0.00881890096296867
"141",-0.023679289444371,-0.037915980237618,-0.0177352428706216,-0.0509649823929915,0.00834255667083683,0.00795993451498767,-0.0229420079317347,-0.0416342608348163,-0.0186846033278145,-0.0106421866674594
"142",-0.019659783009439,-0.0151783461878455,-0.00972217287071175,-0.012954807491945,0.00287217220734992,0.00194408462912277,-0.0276238498937071,-0.0186885671431181,-0.00365571961444877,0.00960418518193684
"143",0.0156432141265879,0.020819946648897,0.0168300081444457,0.032735600191421,-0.00286394645992427,-0.00254636927842233,0.0134942539240877,0.00818594005935203,0.00550363825080957,-0.0114154519572044
"144",-0.0112629458233447,0.00573936175561363,-0.00482708595498915,-0.0204670829573348,0.00723843109824296,0.00413325777753459,-0.0133145835527337,0.0122620161035778,0.000304150842518558,0.00808306373567436
"145",0.00487228413118079,-0.000526991629098084,-0.00762315397038316,-0.00392195424781616,-0.00216370181416514,-0.00277138540805388,0.0156247751151519,-0.00965819512601684,0.002127967743913,-0.00152730162096215
"146",0.00799002883914435,0.00368895972053807,-0.00488840369273658,0.0110559380540383,0.00252369599587499,0.000731587540773182,0.0146852605643852,0.00495875866001194,-0.00060671924768696,0.0015296378393137
"147",-0.0257452002405499,-0.017502348043038,-0.0140350258972289,-0.0431426133852264,0.00664052099120371,0.00645434393420619,-0.0368020461812311,-0.014967222035067,0.0121414935823569,-0.0110728958450327
"148",0.0167594835352765,0.0115793270690636,0.0149466191548104,0.0178469379810804,-0.00727856187366727,-0.00399347376935155,0.0260441796586137,0.00100202051480136,-0.00254918270957627,-0.0138994995789665
"149",0.0106692939639541,0.00255349539514627,-0.00210406080956194,0.00746022956787096,-0.000801214739639233,-0.000121535003467788,0.00404492095975462,0.0158463548225956,-0.000601232739081525,0.00548151681725861
"150",0.0139412752544321,0.0209029717260385,0.00843327619063206,0.033587764477351,-0.012153752785183,-0.00692613149072285,0.0362551177364916,0.0279147526460752,0.00436212375020517,-0.00155763343848836
"151",-0.0296336167007327,-0.0351858606659617,-0.0160282541345611,-0.0413589289883463,0.00139333384257756,0.00562968003498598,-0.00174304204865705,-0.019009535488116,-0.0196195605640062,-0.00780031722738583
"152",-0.00467747047292721,-0.0141774343572669,-0.0141640724595912,-0.0173346238598739,-0.00231892283083512,-0.00146048086103112,-0.03316747097298,-0.00749061640206938,0.0169569357921926,0.00353769611988386
"153",0.00359327168358115,-0.000181149641671596,0.00143666706839629,0.00987862680130247,0.00290487138480189,0.00158348514327078,-0.00416687525129367,-0.0045942888291598,-0.00465672224725844,-0.00705053381947773
"154",-0.0152860912352129,-0.00986056670666635,-0.00286938839774875,-0.0258518992066251,0.00266439904696303,0.00364927252206271,-0.0376565366520808,-0.0214275718173007,0.000452746741540944,0.0031557362828909
"155",-0.0137751893130885,-0.0244859422608917,-0.0165466494370817,-0.0392895837594255,-0.00358107134619046,0.00181861031946884,-0.0108697613782731,-0.0296443649644578,-0.00241369735384378,0.00747162273480795
"156",0.00751575332944476,-0.00290333700256296,0.00219453526144342,-0.0170046983023476,0.010318348829131,0.0038712902887168,0.0257876293879016,-0.0218713888430772,-0.0219264640220684,-0.0171741360556121
"157",0.0183672337648353,0.0186921113611556,-0.00729936110934581,0.0316450816110103,-0.00401662899526656,0.000723475889256031,0.0262820881887806,0.0216510562969028,0.00510207173778587,-0.000794281750049253
"158",-0.00048368943729471,-0.00138274235902813,-0.011029584229626,0.00204525684003798,0.00057604949113288,0.00216801382501575,0.0167014160270376,0.00052109566633729,0.00169206270751987,0.00278215339106791
"159",0.00200506035156067,-0.00277036832946753,0.0126394633876226,-0.00367355068508224,0.00483623249333132,0.00432679616540033,0.0150584095951112,0.0111106507866325,-0.000767859301235019,-0.0015852880109033
"160",0.0118677432613923,0.024722343092118,0.0132161619964117,0.0430152338475154,-0.00160451794752292,-0.0032308657831992,0.00809132598287898,0.0317652141376399,0.00507149223912728,0.00238181403621773
"161",-0.000886291163044617,-0.000813372124453537,0.00724622157358845,0.00510585673089703,0.00344349724006032,0.000359561672545139,-0.00709023768132155,0.00931925099859354,-0.00137620790898463,0.00316823425738266
"162",0.0123530768035416,0.021522884794291,0.00503595697155257,0.0238376141861756,0.00491875591414703,0.000360670206242864,-0.00633235131831067,0.0189612733440492,0.0122493190093194,0.0118436731577627
"163",-0.00930366398071847,-0.00894109873078908,-0.00787392758248906,0.00457984451782001,0.00523632970866483,0.00275926899135959,-0.0135591728296501,-0.00728159206840728,-0.0019663893213373,0.00117050424605614
"164",-0.0219803489199261,-0.024117928171187,-0.00937957082627638,-0.040653430688644,0.00169889353403585,0.00514359079223259,-0.0316153936498208,-0.0221675900915345,-0.00591098790947309,-0.0105221384053501
"165",0.0196216146278609,0.0259039057141224,0.00946838016867857,0.0396040007351059,-0.00271375768830184,-0.00380942675456153,0.026259706831574,0.0218371201124339,0.00731825017949372,0.00945246275909684
"166",-0.00266116478286982,-0.00562120022784751,-0.00649362066835035,-0.00510420059051209,0.00668848397382305,0.00501914510883594,0.00484072652186063,-0.00897267861170081,-0.00408652943847421,0.00195096581230558
"167",0.0098528549158583,0.0171378244547467,0.0217863423266156,0.0258074865956399,0.000787904448104948,0.000238101337688423,0.0199588007870555,0.0139921373222889,0.0109421575558286,0.000389366640277888
"168",0.0100951388998087,0.00961556124986851,-0.00568573219656399,0.0168718484369408,0.000474349598303947,-0.00186146869795278,0.0134954775281559,0.0159091950072008,0.0138305027283752,0.0112884887874316
"169",-0.00865281929561346,-0.0139799537494393,-0.0192994901587937,-0.0151236417006005,0.00801720354138724,0.00621491723255163,-0.0239681720261294,-0.0209334067012434,0.0017793000658568,0.00192459985923144
"170",0.00230069013961542,0.00221518582027569,0.000728928146136898,0.0078272141410034,-0.0025765015897099,-0.00213787584742542,0.00613939174835609,-0.00522274897555408,0.01924220009598,-0.00384172346283407
"171",-0.0139066441039614,-0.0115824266578712,-0.00509846702192485,-0.022559422291246,0.0141508981724416,0.0107153142257608,-0.018712079922633,-0.0164069147534379,0.00769674691117128,0.00655603403984628
"172",-0.00191674350294835,-0.00581461580382225,-0.00878456936550376,0.000756689872971616,0.00775207066079897,0.00223785821895772,-0.0189303515450846,-0.0145120105037594,0.00331465633830019,0.00689651548866221
"173",0.0116600951225811,0.0197051041050946,0.0103399310492716,0.0201887025436069,-0.00076873155247803,-0.00211470345513509,0.0180281958547006,0.018957062850707,0.0129272329965284,0.00228314746503155
"174",0.0025768072695096,0.00326451764431757,-0.00292423711651502,0.00355822391063598,-0.00373887135706752,-0.00247429696926615,0.00179854073470564,0.0101329952503719,-0.000850794137158162,0.0106301868737808
"175",0.00703290221928121,0.00562882648844099,-0.0073313124260922,0.0110784259223735,-0.00894145572306715,-0.00590328742054691,0.0183676815985205,0.00970233910337681,-0.00539308835357777,-0.0075131534517725
"176",-0.0000670514595694227,-0.009970379264155,0.00295422386308197,0.00197171808535712,0.00144746137067209,0.00130680548090023,0.00474617254205034,-0.00716644733417116,-0.00128430361631549,0.000757043374380428
"177",-0.00537279791631484,-0.0167839579007155,-0.00515469201709218,-0.00634225233858421,0.00478252230673282,0.000592388221638096,-0.00188940442077123,-0.0247700015832637,0.0140020435491368,0.0117245866427997
"178",0.0294397529762471,0.0420484269914554,0.0103628920705598,0.0484228617669347,-0.00752697611800202,-0.00106612870723555,0.0311020946383482,0.027754310310224,0.0102859798466115,0.00373824050057459
"179",0.00590296447276772,0.00353475156768801,0.0109889323144736,0.00454816181436701,-0.00925743077078622,-0.00356099074511107,0.0203278018419573,0.0193127761469973,-0.00376564869312324,0.0085661949880711
"180",-0.00704192207032606,0.00223399125260837,-0.00362335574655792,-0.00313459336338662,-0.0189117201248198,-0.0113144202784702,-0.0122108296059477,-0.00851018409565873,0.0180596528069437,0.0155096524025742
"181",0.00269861135894489,0.00642953517601641,0.00218176733748243,0.0132774657815591,0.00848981169105945,0.00505940017618944,0.000260119668365366,0.0131568700741951,-0.00522559123727184,0.00690905679580123
"182",-0.00184253499098197,-0.00170352287660636,0.00362854849763972,0.0124138532757738,0.00284518501920572,0.00131851266018912,0.00858593300292965,-0.00145187249113188,-0.000829375218654893,-0.00180574604944927
"183",-0.0019777340877507,-0.00392505779696128,0.00578448758991312,-0.00374655844856675,-0.00351698982310356,0.000120221214905847,-0.0165534175425976,0.00226160943029763,0.000691795803704931,-0.0072358181019565
"184",0.00528447480960259,0.00436874230940432,0.00862686273558522,0.0133333429986002,0.000910541507065155,0.000358915230032952,0.00569022194158708,0.0169250447707769,-0.00456244975632647,0.00145768792851686
"185",0.00591344315019837,0.0119403259719932,0.0228085107054081,0.0148448482260353,0.00693921651111085,0.00322978282897712,0.00947341546171621,0.0112536391858253,0.0097221805555554,0.0262008927706412
"186",-0.00333144175767919,0.00463540350239167,-0.000696947654528324,-0.00631664958041123,0.00225903763483948,0.000357958107760181,-0.00325845910770994,0.00705288403263893,0.011141747364859,-0.00319145367419116
"187",0.0112724918214766,0.0100671701802122,0.0111572895218768,0.031448666523163,0.00571437607761416,0.00119662068804582,0.0265462942119317,0.00498086652666285,0.00530540048142014,-0.0103167347210077
"188",-0.00136039398524035,-0.00299006219371301,-0.00275857099333698,0.00681168204821292,0.00315037016741315,0.00215103625394319,0.00917227598582504,-0.00263262852442792,-0.020974343140072,-0.0201293040553866
"189",-0.00201212439030607,-0.0036653775609492,0.000691709834153453,-0.0302839006581719,-0.0029164908554592,-0.000715304892912272,-0.000252296620582459,0.00155242407057021,-0.00621970991623244,0.00110047505025279
"190",0.00156103054322698,0.00526765961410125,-0.000691231702387274,0.00996708927285206,0.00382524841282961,0.00178951786947712,0.000378583128679111,-0.00465110074952335,0.0134909731991384,0.013924485602435
"191",0.0118813321572453,0.0075687015309307,0.0131398090156567,0.0333551754333259,-0.0107577605500545,-0.00881568404042121,0.0198155035809673,0.00934579294627991,0.0072732122708985,0.0028913363212475
"192",-0.00532572639043827,-0.0114743748371521,-0.00546063061845636,-0.0106320642025607,-0.000793607052438472,0.00360617295635191,-0.0111382890219468,-0.00925925783967396,-0.0118529015843896,-0.0209009532259744
"193",0.0094179991421186,0.0125261341712128,-0.00274538023614357,0.0155724964476918,-0.00124609461681624,-0.00311420482962688,0.00575694864963139,0.0171339537348463,0.00772090180230101,0.00699301195640767
"194",-0.00166115870147709,0.000412289764066376,-0.00206496266409273,0.00133069117470463,0.000567020233888327,0.000962095610222757,-0.00136899841642946,-0.00137779149213157,0.00369414440794325,0.0116958755188288
"195",-0.00480140800402573,0.00412211510530236,0.00137960340693843,-0.00879541404485895,-0.00102075929197709,0.000119405195059707,-0.00672862455176271,-0.003987335471755,0.00749731451066915,0.0111994302013048
"196",0.00553220629529116,0.00615777720513466,0,0.0182580632466007,-0.00488289973266787,-0.00335989686195093,-0.0072766514477911,0.000769761450125195,0.00920027010146018,0.00464463410506832
"197",-0.0084443244571738,-0.0087314557649053,-0.0117078910424115,-0.0122254448913971,0.000227626326071428,0.000962849986003489,-0.0205990056725133,-0.00846171902843795,0.00737368319472775,0.0170696735864164
"198",-0.00793470539053998,-0.0113596932094249,-0.0181187116182485,-0.0185339440601711,0.000342863427091666,0.0027674065335006,-0.0166452240497506,-0.0217223544621982,-0.000266116585921239,0.00104887679717081
"199",0.0030563534045791,0.0122396513572509,0.00141948607458908,0.0230870835848402,0.010948776209369,0.00611806233140566,-0.00275534241778697,0.00475847482491232,-0.00825350073535003,-0.00523930066369616
"200",-0.00363008495480188,-0.000493341667171521,0.00425237841036519,0.00505716369100706,0.00552748226758082,0.00381502919895493,0.00263141778472264,-0.00552476553110881,0.0201342281879195,0.0179073168434274
"201",-0.0261568307025725,-0.0198337454580347,-0.0197598689063124,-0.0427674747376316,0.0149218181924371,0.00855272044634603,-0.0322832010645902,-0.027301964609576,-0.00394740789473691,-0.00275953735000611
"202",0.00581265261813013,-0.00503799983534658,0.00575925589957116,0.00722736825637726,0.000111249906017852,-0.00188443169151697,0.012340438010199,-0.000489445835774038,-0.0145310309589576,-0.00276717346854638
"203",0.00810429694177284,0.0156118292291763,0.00286344637619873,0.0277237337641281,-0.00132657907110234,-0.000236117444040507,0.008707345910973,0.0179588551928092,0.00844510746501625,-0.00693725997684724
"204",-0.001845411609804,-0.00124621882870557,-0.00428288375823849,-0.00653765220475822,0.00741582160885135,0.00507409191497921,-0.00398429148804946,-0.000160040765461389,0.00385476523243011,0.00349284216203993
"205",0.00237700457054557,0.00582360284993011,-0.00358415343191221,0.0127138836447285,-0.00340635543008172,-0.000821191158103085,-0.00266659429152161,0.0131539059942438,0.0067532047174208,0.0233204754837524
"206",0.0117224899154966,0.0168732558813505,0.0172662266236352,0.0283262214226896,-0.00231458151301311,-0.00246864553607629,0.014706069819606,0.0186825632220284,0.0218335265268121,0.0153063169226604
"207",0.0033203990884072,0.00618216907562319,0.013436997709191,0.0230063673621512,0.00386738064513459,0.000824993308214284,-0.00724654580945172,0.00326394644570782,0.00553483059506155,0.0164152409450689
"208",-0.00694264236790387,-0.0072758579543809,-0.00488473599296724,-0.018890642352529,-0.000550361495205709,0.00105923233175353,0.00451231473509139,-0.00325332775813503,-0.00985669444994774,-0.0224126033472398
"209",0.0103881918854678,0.0146580010603905,0.00701253751548214,0.0219437202299815,-0.00903060561374913,-0.00670275325489977,0.017967756457872,0.0219147336994612,0.016418940308182,0.0283210275855652
"210",-0.0234076406180154,-0.0244780356450192,-0.0125349330683192,-0.0403733972485415,0.0129928676373643,0.00816154937166158,-0.0356907933063755,-0.026768181289057,-0.00877643059871147,-0.0127869289061899
"211",0.00112535934169955,0.00822697432600195,-0.00282073673428684,0.00567200865125583,0.0031956069879111,0.00271092839574072,-0.0197844597118804,-0.0078137199719136,0.0243808802771717,0.0215875633978628
"212",-0.00760521999713937,-0.0134640286649623,-0.016973164125327,-0.034769259994161,-0.000439451863856077,-0.00117470865264402,-0.0142796734087554,-0.0195305948681092,-0.00100215455337194,-0.00650202454672566
"213",0.0134618332236813,0.0140612661179207,0.0115109577718935,0.0379479042607913,-0.00483543235052142,-0.00176567942143424,0.0104470484016754,0.00883533995538044,0.0210658307210032,0.0261779946862162
"214",-0.0273559572831849,-0.016068569031905,-0.0184921865848976,-0.0318586744011286,0.00176670235450294,0.00365396189781153,-0.0337751102876964,-0.019586256263014,0.00994716934790607,-0.00510201048791581
"215",-0.0050706899647025,0.00887005698693821,-0.0159420927589582,0.00511161900718893,-0.00176358662186582,0.00223061538501579,0.00627817827468502,-0.0035727948149521,-0.000121534536029588,-0.00256400139839019
"216",-0.0137262724771599,-0.0230073248121018,-0.0132549061654967,-0.0235219965966874,0.00850321637640827,0.00597687803977909,-0.00340295834903925,-0.0203749252337623,-0.000608087050659512,-0.0003214058130524
"217",-0.00992156258815913,-0.0159799210568442,0.000746243634889732,-0.055338608770199,0.00361294948962598,0.00174713760759238,0.000142583761104875,-0.0257904095710222,-0.047213397420297,-0.0218579729895122
"218",0.0304801197385598,0.0286324291648321,0.0171514465916318,0.070640964289437,-0.0037091914366828,-0.005115918508942,0.0358463104616982,0.0401366964163938,0.0104725411057773,-0.0190600112852922
"219",-0.00276877381441232,-0.00290788554751431,0.00293281335819273,0.000965440041944765,0.00109479346469188,0.000701452458945262,-0.0146938966173247,-0.010673199746856,0.0146612229021277,0.0224454312693505
"220",-0.0144241498350719,-0.0166670055567286,-0.00877214973930718,-0.0230221350201815,0.00940723690721712,0.00560584368622519,-0.00557475992030665,-0.0182571906366428,-0.0290234433112039,-0.00982962716745794
"221",0.00171796023925008,0.00423731845688913,-0.00737490466435464,0.0123747751532897,0.00140854852807015,0,-0.0190610287544479,-0.00422667563616963,-0.00256570888642882,0.00330906930670882
"222",-0.0139243049929322,-0.0270040416028392,-0.0170874628649808,-0.0460988183844845,0.00649341792972358,0.00720091395911893,-0.0191455772453463,-0.0280135766728004,-0.00655951125401932,0.00758579294261863
"223",0.00612141915924025,0.0222895690639009,0.0264551379273028,0.0274692790548057,-0.00107478988771115,-0.0026519509811066,-0.0233066015090455,0.0155462578315058,0.0288710908563203,0.0248772327886559
"224",-0.0204643933183575,-0.0184947296327678,-0.0176732459370562,-0.0503517530816783,0.00581124154859824,0.00786164419439239,-0.00745719330342809,-0.0223603201521001,-0.00138417010967451,0.00127765068033292
"225",0.0172923383039558,0.0215226339981829,0.0224888787853839,0.0295494746945355,0.0029967844923553,-0.00298205760680004,0.0190835596031045,0.0362421913556661,0.0238155112926473,0.00925023354463761
"226",-0.0220632962603908,-0.0197156003663693,0,-0.0396934217180184,0.0197371564880777,0.0136914564984105,-0.0376000710963001,-0.0290325288115001,0.000615421538461502,-0.0123260774232595
"227",0.0114930446899757,0.0125162064953597,0.0161290991221612,0.0382957741172469,-0.00952137395792396,-0.00930713556630525,0.00735444866462553,0.0307747592198213,-0.014760208557434,-0.00800003976861519
"228",0.0319845925459554,0.0323956331829625,0.00937937127226163,0.05478083510984,-0.00675940609971037,-0.00355181117985592,0.0468440896748827,0.0154369513809964,-0.00661670428506134,-0.0122580734124823
"229",0.000339768860850409,-0.00908317331194908,0.00357423512286581,-0.0122582736469384,0.00861436084556422,0.00563430587923808,0.00799078934912489,0.00133637178115231,-0.016212152821415,0.00228622915887211
"230",0.0100555848153883,0.00374991035272743,0.00213637357966712,0.00849135184401817,-0.00485083278549669,0.00137196146392027,0.00922392128004268,0.0060063102224257,-0.0122636562629492,-0.0123820652419223
"231",-0.00659266844074091,-0.00356992476656159,0.00142161324348478,-0.00867879222144252,0.00793588254949995,0.00395184599084697,-0.00728300985487573,0.00364817255104222,0.0124159208484222,0.00725844226775885
"232",-0.00893800134457723,-0.00599898234746155,-0.0106458620198988,-0.00261372577751451,-0.000105574048168577,0.000913571513384337,-0.026183525054548,-0.0133840751440543,0.0143076522011707,0.00458558632946859
"233",0.016739684437155,0.00813030574084483,0.0186516198118354,0.0444128423259196,-0.0119273191205331,-0.00376258010154951,0.0285124041974743,0.0217719617400531,-0.00969779572549634,-0.00749915544072055
"234",0.0143134583420981,0.010643282100893,0.0126759313644227,0.0157424072528416,-0.00875939720701124,-0.00526444513974844,0.035909550407744,0.0136044095319876,0.00941124288736761,0.0180682734706157
"235",-0.000198411226577488,-0.00255062359784053,-0.00904037163438642,-0.0118554090044461,-0.0112082541641623,-0.00644191806142425,-0.00485346276338294,0.00258700659191069,-0.00970146114269388,-0.00322681525340973
"236",0.00775257923736294,0.011217481575738,0.00280694479509891,0.00031232023460448,-0.00599529709538726,-0.00231689334277208,0.0250804705043406,0.00403248265779599,0.0178117307331229,-0.000647459196076228
"237",-0.0274196304252033,-0.0268354833338015,-0.0216934097981948,-0.0423538252397522,0.0196278366064271,0.0136953088301053,-0.0572244264867664,-0.0224903073603734,-0.01450005,0.00874629264896143
"238",0.00987125934247923,0.0233846155706041,0.00786829479934426,0.0300066451084842,-0.0103242670560819,-0.00835715470961051,0.00317185730139968,0,0.0209284891389392,0.0272961382131933
"239",-0.00207557521876489,-0.0197378104944859,-0.0205817847059131,-0.0274859022823994,-0.0108660778206022,-0.00739002074205919,-0.0172467588081597,-0.0164331059277806,-0.0247235439116299,-0.0106282956909713
"240",-0.0126796451593891,-0.0252318538871114,-0.0391305629749911,-0.0238343528014023,-0.00461331756283867,-0.00290818490082179,-0.0302715613402386,-0.0342525768703734,0.000254738853503245,-0.00695106564738879
"241",-0.01426926331261,-0.0173996326749936,-0.0173454661325906,-0.0426281805627159,0.0089394507707492,0.00595035380915854,-0.018097134481844,-0.0501731684652021,-0.0049668876069876,-0.00489079563714301
"242",0.00558387149317108,0.0109910612815065,0.017651642092694,0.0274539731013916,0.00645331848524822,0.00197102726198173,0.0129012609219512,0.00273195060093023,0.0143351215026926,-0.00425944207669848
"243",0,-0.0101812135081012,-0.00678726461657231,0.00651120057195853,0.0132600434821057,0.0079852003735672,0.00833964157206601,0.00999153274618991,-0.000126208201892797,0.00954259968372395
"244",0.00630655214186171,0.0039226842720208,0.00379649613974276,0.0054577786700325,-0.00214543359348196,-0.00160610758815205,0.00375963915843647,-0.0062952114866569,-0.00719333688019519,-0.00423733058600284
"245",0.0144151609778256,0.0145869754090144,0.0151284328503842,0.0301568821923941,-0.01461881777527,-0.0072459305306537,0.017078338731487,0.0130323695503434,0.0181771963436428,0.0117839818799261
"246",0.00742607720432775,0.00679761266296208,-0.00165607939764778,0.0169132347786316,-0.00469040330589365,-0.0028967692742452,0.0272503547478133,0.0189192180827122,0.000499388277138246,0.00744093606279606
"247",0.00214432934521569,0.00550276233892943,0.00452499824469776,0.00518334426279243,-0.00876827810216574,-0.0047626570949092,-0.0166331816219517,0.0150307645577412,0.0172198404943829,0.011881835103565
"248",-0.012571187990667,-0.00277987689406922,-0.0157660150402722,-0.0230761278522646,0.0109015968001049,0.00671321622732979,-0.0194546744041096,-0.0243899860432898,0.000490689419431423,0.0034910490379898
"249",-0.00250587550955694,0.00836241993013087,0.0114417916288641,0.00376108874281167,0.0155934663191817,0.00803099241763006,-0.0147414815211305,0.0157143024013324,0.0176557385398661,-0.00316255885803629
"250",-0.00739960797394079,-0.0122669113543042,0.00226224680840637,-0.0120290096388749,0.00605600313901156,0.00461829564975291,0.00305371744441496,0.00123034978734649,-0.00650603614457834,0.00126896397825904
"251",-0.00875443213513682,-0.00271103863760136,-0.00451460160058648,-0.0165006210589274,0.0144023564329676,0.00712544073061117,-0.00837153985290651,-0.0043898632550694,0.0291050452231998,0.0275666024282257
"252",-0.000483197740811514,0.00175380025531746,0.00377926803309614,0.00899761447492531,-0.00137709450501189,0.00205431529570577,-0.0323869156057448,-0.00370356753840073,0.00836670977649412,0.00770883958221713
"253",-0.0245064505079465,-0.0234611774522098,-0.0256024938350035,-0.0300368890857619,0.000210938072806366,0.00262018786786533,-0.0317258521213297,-0.0219506570349396,-0.00514202407385755,-0.00581387407030654
"254",-0.000849014498128575,0.00502016031093167,-0.00618234577647636,0.00732711082994064,0.00434951173741882,0.0018160813225756,0.00933833520252647,-0.0162897587377726,-0.00422882664967084,-0.0181595601336975
"255",-0.0161483294004671,-0.00909840705034792,-0.00233268359840499,-0.00775401648514273,-0.00116147123742305,0.00215468993223067,-0.0363580434001537,-0.0220791884382113,0.0237112430238733,0.00909093024415042
"256",0.0105100787933279,0.00414099936058232,0.0218237725612547,0.0327800947462984,0.00190318687810231,-0.00158450839249835,0.0197071882646258,0.00564459743542045,-0.00265033420892291,-0.00994093566611409
"257",0.00655422285641283,0.000806632649623884,-0.00839044767382313,0.0117849340841945,-0.0135091543699712,-0.00271956384394434,0.0132145740922223,0.00187104532115012,0.0196417901915036,-0.00470664262171938
"258",-0.0080686298979129,-0.0173773854334711,-0.0169232602787455,-0.0281268934915615,0.00781019587872489,0.00636271815805789,-0.00163025789164839,-0.0252099891132497,0.0037393994334276,0.00914241888765055
"259",0.00806281352481197,0.0165909001059943,0.0125195634913327,0.0147085669599478,0.00371546558109581,0.000452260940307037,-0.00277648251352303,0.0153253247211822,0.0108376493376012,0.0124962089895626
"260",-0.022013047442261,-0.0312949336084282,-0.0278207675380027,-0.0452317931932623,0.01121117417513,0.00654600295452901,-0.0260354415815468,-0.030943294128266,-0.0173107324401304,-0.0123419810154484
"261",-0.00861222294791897,-0.0216603844947462,-0.0182827188441834,-0.0416108779040313,-0.00721712223338911,-0.0019063267251539,0.0129452808266239,0.00272555127984253,-0.0146607686023587,-0.00937191995711351
"262",-0.0259167944548944,-0.0142874542889451,-0.0137652995420589,-0.0291162431415638,0.0129586958333872,0.00808752442221761,-0.0121159967875764,-0.0108736043301751,-0.002306770552714,-0.0129297788189532
"263",-0.0102672655339821,0.0010562309951474,0.026272653813346,0.022813333449303,-0.00686446648949468,-0.00144782893675777,-0.00840071036880452,0.00706708724023963,0.0106358150289019,0.00383388391305206
"264",-0.0101465445653797,-0.0312590475164453,-0.0368002996564093,-0.0251110659297117,0.0106815065598362,0.0111592404519218,0.0337176050889958,-0.0183234736199698,0.00857927267397107,-0.00350091581404965
"265",0.0240205095651824,-0.006532805513361,0.00332234213955074,0.00636341590498901,-0.00227900071582676,-0.00463570461119889,0.0817898812090188,0.0127084896413487,-0.00317567206931324,-0.0188438187034397
"266",0.00844182481259237,0.0297897453072662,0.0165564518811327,0.0194220031928309,-0.0200442864303627,-0.00909135990734145,-0.0195455141035777,0.0284313842903927,0.0249175449416035,0.0247395512072714
"267",-0.0144456623759296,-0.0201240723173385,0.0154723487868418,-0.0152117216836164,0.0168502328815257,0.00928740203435363,-0.0139080580513887,0.028599197606576,0.00244228458165452,0.0222363674138357
"268",0.0165366759089565,0.0156993102035239,-0.00561341590425157,0.0247447780155516,-0.00375175160241659,-0.00365962480155058,0.0371413703287975,-0.00185428823784717,0.0160575520689628,0.00466139951663203
"269",0.00495375796357345,0.00767954360867651,0.0169352881377509,-0.00490240327090907,-0.00679953996276295,-0.00400448222162986,-0.00604427667667284,0.00185773301031733,-0.00653948773841961,0.0083512203980638
"270",-0.00735742783810067,-0.00347290595089489,-0.00475815019849912,-0.013162729067685,-0.00653009789639025,-0.000447058271186074,-0.0234112342498558,-0.0157562276004234,0.00998349950667032,-0.00858889055647272
"271",0.0182340314955101,0.00948687159628148,0.0135458384965639,0.0200448129448243,0.00710269201828662,0.00514109236266402,0.0238171310083484,0.0169496676109782,-0.00716919415966089,0.0049505395663092
"272",0.0160879552107447,0.0138090597709453,0.00864796576479931,0.0199427276214548,0.00601152197229782,0.00324523852716418,0.0389236866984439,0.0203704115191787,-0.0224289272991482,-0.0175493094837592
"273",-0.0126091681466669,-0.00813454019122584,-0.00311793579152186,0.00308007378271524,-0.0102920108552332,-0.00555890569249184,-0.0155133948008984,-0.00381146851172398,-0.00279798551310539,0.0175493516543039
"274",-0.0267740067158313,-0.0500669277514108,-0.0336201876603119,-0.0538380223247271,0.00764045268664026,0.00704396553576991,-0.0316633909446961,-0.0435418933961362,-0.0159371271815292,-0.00831537447744168
"275",-0.00805189214374791,0.0055215984166781,-0.0129445951101625,-0.0163763112482448,-0.00305445899545742,-0.0017755240341929,-0.0191893719896009,0,0.0144844548357663,-0.00465840677163776
"276",0.00661378819324954,-0.0108827311449352,0.00573744778571483,0.0169558841782369,-0.0215457131079042,-0.0112337842191786,0.0241041760539755,-0.00857127577429617,0.0101180554283773,0.0121684457745848
"277",-0.00642103209191092,-0.00353267970778981,-0.0252646615301564,-0.00188633017367545,0.0114417183567666,0.00843508627623901,-0.0310256591101195,0.00192148525309954,0.0127991321713774,0.0299014221653737
"278",0.00511008387172107,0.000911821031994497,0.0100332861921568,0.0123961825026566,0.00416301098492555,0.00223200808275736,-0.0200315800254692,0,0.00362639560439559,0.00658490632753428
"279",0.00927112619522297,0.0254022211461165,0.0149006808018453,0.0161266228889894,-0.00595217716925289,-0.00211468387435776,0.0315464744600713,0.0134230903585739,-0.0218986089587516,-0.0202200517606466
"280",0.0102228545362462,0.0141133648542773,-0.00734090555399625,0.0224835735220013,-0.0105850491233218,-0.00423866079038626,0.0046811033088523,0.00851458115311976,0.00123138920337218,0.00819414455935585
"281",-0.00879967906669832,-0.00778587917254048,0.00986033226559879,-0.0128629998182513,-0.0146967979683866,-0.00548817864988549,-0.00745442181663181,-0.00093815527673069,0.00301874993249651,0.0201685945015921
"282",-0.00022193589834385,-0.00392301409333462,0.0122050012364106,0.00713427358413532,0.00767797513215163,0.00214038505614189,-0.00406827473010085,-0.00187825747967396,-0.00624230304583995,-0.00472116848927839
"283",0.00281179607841464,0.0125058962501865,0.00964651765888513,0.0130827302418146,-0.0101218461076743,-0.00719245144346414,-0.0174393901083244,0.0169329767629849,0.0272574306840732,0.0326120194826895
"284",0.00295174902473239,-0.000486494024286244,-0.0207011714685306,0.00834780442100302,0.00692677724257584,-0.000906144951648313,0.0233452357357713,-0.0129507650824301,0.0181261843606424,0.00516786232688937
"285",-0.0083137469206912,-0.00136185034312186,0.00731743063966306,-0.0140100388687558,0.0105917452414352,0.0103112259363585,-0.0226561573709664,-0.00674802827200005,0.000107271559572464,-0.00542700647917216
"286",0.00615787716821914,0.00964630939727806,0.00807127462397017,0.0134195085297415,-0.00572663487032488,-0.00280448417950141,0.023501422856975,0.00490706858220835,0.0015013297587132,0.0137852753837973
"287",0.0126090102453824,0.0147653744059544,0.0208164347615836,0.018623240047525,-0.0102149451960506,-0.00663540288876963,0.0309275804360569,0.0140844335623445,-0.0069600707459051,0.0096317030604518
"288",0.00750007689531462,0.0194958962902108,0.0109805452975136,0.0132080919192838,0.000329202214973678,0.00249105509561209,-0.000606111530903508,0.013888890409165,0.0104593597252396,0.0213242670851113
"289",-0.0010119842506715,-0.00335844015960285,-0.00543077102479461,0.00843907175955994,0.000877972425131546,0.00237143994022904,-0.00712540753755186,0.0100457903383904,0.0114182052226892,-0.00137369983327418
"290",-0.00976699816465776,-0.00393128314035807,-0.0109203050166514,-0.0107495669808851,0.0177648024310801,0.011716991699084,-0.0207666137554956,-0.00542546061920868,0.0127663959988014,0.0096287237141659
"291",-0.0222840364918048,-0.0247130624247834,-0.0118296337203617,-0.0397525375660617,0.0153011010639159,0.0106902255310655,-0.0174644551881402,-0.0334541138039408,0.00197939372808409,-0.0163487644500253
"292",-0.00239133693885185,0,-0.0007982014143042,0.00544360079109474,-0.00257851125283426,-0.00254215723564521,0.00539607714480983,0.00169300826023022,0.0110209814930338,0.0146813734667879
"293",-0.00382015543469827,-0.0112727219654277,-0.0231630528085012,-0.0232226916846783,-0.00971798579815875,-0.00376652258883048,-0.00805054174293507,-0.0159628390441048,-0.0211846775233376,-0.0035489822077398
"294",0.00631605924380585,0.0109141448362351,0.00572337527661637,0.0210033259973603,-0.0119699411510422,-0.00433773645179603,-0.000954965747412939,0.0160308482455345,0.0266862891363731,0.0219177486587276
"295",-0.0206976005616776,-0.0113750687645028,-0.00894272130685181,-0.0342854905399719,0.00534808790919006,0.00804293314164073,-0.0458747705348299,-0.015965394754294,-0.0124846601260268,0.00750686883795959
"296",-0.0103009596979171,-0.00887236371943712,-0.0147661192760029,-0.0138319673747022,0.00130270712304847,0.00343506068195731,0.0100172045749469,-0.0112622497391703,-0.00424874611398962,-0.0101118449885799
"297",-0.0131832105447911,-0.0102315181472908,-0.00416319904356666,-0.0175499718582049,0.0147450679627616,0.00717823241510462,-0.0161985725944093,-0.0173743233014056,-0.00228944748837334,0.0188172265118327
"298",0.03593786233327,0.0318060916567073,0.0292641498105235,0.0672569197708202,-0.00854707873999028,-0.010855595110182,0.0710682192519245,0.0451867719598,0.00125164281052537,0.0155672258795234
"299",-0.00935146192180358,0.00250440415903164,0,-0.01852633504349,0.0192904546327071,0.0115293035958108,-0.0214895318743102,-0.0203007926185373,0.0106261487785426,0.0109120036113952
"300",0.00220782569107514,0.00490075551393998,0.00324957017689176,-0.0091099438037513,-0.00782348889415729,-0.00526055845817619,0.0125034199044645,-0.00230195961050184,0.0137098646797265,0.00102792855388745
"301",-0.0154960459555179,-0.0253393237489293,-0.0663968447882647,-0.0354517642378482,0.0123611285678438,0.0103557674066883,-0.0163075102992037,-0.00576950328543779,0.00376248744203722,-0.00128365835410771
"302",-0.0101071171840292,-0.0171689341874067,0.028620983920514,-0.0247066080866766,0.00768384218579565,0.00501580148824887,-0.00675980701038559,-0.0348163773177921,0.00466010540634287,-0.0401027999348437
"303",0.0415430896640618,0.0303454485724159,0.0286678071977582,0.0519937515595033,-0.00386504871149074,-0.00683535235876531,0.0510449787702609,0.0320640107524293,-0.0269234451330734,0.0222280619906789
"304",-0.0247696560838003,-0.0382678071647257,-0.0303276458464203,-0.0600520154488141,0.0165689270687448,0.00863062997236153,-0.0109467622055005,-0.0194172298379762,-0.0358549119170984,-0.0432275970356528
"305",0.0185227943093058,0.0126927967412982,0.0185964974075654,0.0168423485573259,0.00247604999235751,0.00216585216163989,0.041777003596891,0.00406240140074687,-0.0336414119342067,-0.0402519045767038
"306",0.0199877734052689,0.0179052901480585,0.0307054477518849,0.0383356393047503,-0.0193452868392384,-0.0176157607581,0.0170581680378861,0.0392700655161671,0.00211315750803442,0.0182596148216252
"307",0.000964799234028479,0.0177853737606517,0.0104668310480676,0.0153523543127658,0.00419710471752666,0.00352072996003283,0.00788446508107032,0.00954207934766793,0.0291898452650354,0.0100869355330777
"308",-0.012235387945058,0.00384045511313658,-0.00796827715028392,-0.00811339236729092,-0.00417956265538855,0.000766725750176001,-0.0264201940627258,-0.00378080732059993,0.0115388759342541,0.0299583839720059
"309",-0.00315342579205946,0.00124389864929397,-0.0032126630495819,-0.00483317884915191,-0.00703086942291509,-0.00131458965034981,-0.00424514520048536,0,-0.00362477600347211,0.011042175200366
"310",-0.00956449794773873,-0.00487230672132932,0.00402901085848462,-0.00179381181273353,0.00972167747785324,0.00394885717336946,-0.0153777401818236,-0.0153700382196028,-0.0169056496565979,-0.0237079151963853
"311",0.00349766878885216,0.00806367122116169,-0.00722297594625354,0.00591404672286111,0.00355885281275592,0.00174819007520344,0.00664915964963564,0.018500847658026,-0.0159990536351454,-0.0240109860613007
"312",0.0351593072162013,0.0318066362195559,0.0291025993673668,0.0383986057201606,-0.016274819852682,-0.00874346491225375,0.0491552368848565,0.0454119779377657,-0.0392655994130915,-0.00559131338682139
"313",0.000659127698401152,0.000369007484574135,-0.00157103522725277,0.00071654064810267,0.00212841708543787,-0.00331232345506616,0.00424622042625811,-0.00271550004147103,0.0277457514650501,0.0298003766841444
"314",0.00248673369260111,0.00166083847926246,0.00472071322948597,0.0121743290493093,0.00223191468944717,0,0.0204110551620138,-0.0018151560355405,0.00168030699048871,0.0054601548488511
"315",-0.00109436727174517,0.00543393224295374,0.000782914136891355,-0.0040329336084548,0.00911560243425802,0.00764355704414732,-0.0162881870624639,0.000909709303385853,0.00928206238608942,0.00705930535222699
"316",0.000511708991401516,0.00494704885317243,0.00704221430281904,0.0132839202663499,-0.00525191760294497,-0.00659680272691143,-0.00232393979699963,0.00999076739391747,0.0101938836565099,0.0107847322711923
"317",-0.00102232868343444,-0.00911573944499544,-0.0147628622245666,-0.00546823674552899,-0.00348368488326212,0.000111103063239026,-0.0125197373436509,-0.0151081267410563,-0.0089941868815222,0.00400083423797892
"318",-0.00723589446850081,-0.00386371764772708,-0.0149840939721547,-0.0155784288570125,0.0103831215540833,0.00597545843642133,-0.0203454440166493,-0.0189917700803127,0.0214720868062444,0.0167376768781422
"319",0.00139889786225433,-0.0029554807352794,-0.00320298174149425,0.0143211044137508,-0.00335548326572432,-0.00396031462273139,-0.00210648639204125,-0.0087490282423518,-0.00563445654313077,-0.0044422060963667
"320",-0.0194090197575291,-0.0163022718032189,0.00642601013829025,-0.0163073109389673,0.00673485254241091,0.00430654413464859,-0.00361968605473484,-0.0101412848178378,-0.00512143418725408,-0.00393697157603001
"321",-0.00337401362878886,0.00197733570370562,-0.00638498019085121,-0.00236869248263982,-0.00585339000454099,-0.00252841213729593,-0.00544861570235577,-0.00986516432957951,-0.00208107331606555,0.00685105097014449
"322",0.00233247286414495,0.00488691932724628,0.00722904764334942,0.0117259766111306,-0.0124069044886721,-0.00451951415455032,0.00517428682845367,0.0136043205818777,0.00603669184461975,0.0120387266780331
"323",0.0270937846017274,0.0301131708342173,0.0318979685291314,0.0295786522312789,-0.00979487263689172,-0.00675518662293229,0.043149097449859,0.0302455697037949,0.0175648366762018,0.00956836643833903
"324",0.00146156558511512,-0.0128008209788623,-0.0146831182288778,-0.00725116400546122,-0.00172031574241849,-0.00234057169263169,0.00580558560992639,-0.00422007683435854,-0.00761229787538231,-0.00461070342382686
"325",0.0104339915922638,0.0121388990567661,0.0274510173442382,0.0150957180906437,-0.000861344661322483,-0.00100557505829491,0.00101052403802604,0.0068176983117505,-0.0209593241348168,0.000514571753596815
"326",0.00050548847977927,0.00254422217806161,-0.003053325016102,0.00507098068476797,0.00398810680155703,0.000111620283384628,-0.00994697090209695,0.00311169702192582,-0.00408301685887158,0.00128607698844219
"327",-0.00440281475766535,-0.00879120698549285,-0.0191425423767695,-0.00927308757041378,0.00343606200400481,0.000783019921675399,-0.00465928732774068,-0.00437875754081818,0.000221573407202191,0.00616493979980648
"328",-0.00159483459042287,0.00128039073013797,0.0109290901965728,0.0143840917962419,-0.00331701771497839,-0.00100558281114049,0.0115561158919444,0.00293175893868014,-0.0116317274276636,-0.00944611904816373
"329",0.00435693248152624,-0.00392670712821319,-0.00772208072126779,-0.0128228419749586,-0.00848093631823921,-0.00783175397642144,0.022993675052934,-0.00877042570112285,-0.0224164982916779,-0.0167525302708712
"330",0.00925373543829422,0.00980939541551895,0.0194552134077282,0.00735360180449662,-0.00584630401237418,-0.00135325874136127,0.00339300845893242,0.00460817793402879,0.000573217145457328,0.0183485356086419
"331",0.000215028050339239,0.000726061013337942,0.0183203680168176,-0.001910222151007,0.00304916681223544,0.00180717762782501,0.00225375887106538,0.00642221553818123,0.00481270785422394,0.00231666710798772
"332",-0.00393913787709688,-0.00816475389299465,-0.00899515723952016,-0.017704538299968,0.00380030325596814,0.00180367645271073,-0.0144782985612923,0.00182300046724282,-0.0214392058059254,-0.0241397522296555
"333",-0.0058959503750754,0.00301852211712728,0.0045384827863435,0.0205982590036988,0.00713849914198939,0.00314961862061836,-0.0175442712067534,0.00873542055371668,0.00978911571586338,-0.00184207728080377
"334",0.0206858528088727,0.00729548054938989,0.00903600184791276,0.010637072355745,0.000065325429514651,-0.000112613173389398,0.0235194642986001,0.00739702265578979,-0.0306982566486265,-0.0232005671045774
"335",0.00276317781265245,0.00153893335390576,-0.00223852124587542,0.00958037585484983,-0.0126110630352317,-0.00810135127026612,0.00170205686188551,0.0109232603845866,0.00702469358315727,0.0253710588069842
"336",-0.00480468331181227,0.000632639442437632,0.00149574114155548,-0.000735199974755796,0,0.00147527783693513,-0.00240685753453329,0.00212603418876212,0.0199810234102384,0.0207949517827233
"337",0.00866278103766205,0.00505870821428922,0.00448063529868348,0.0111683642098379,-0.00720373512556605,-0.00317154663207353,0.00794866059100086,0.00212124669140712,0.00417294554907666,0.013151143431118
"338",-0.01781065787812,-0.0171669046866697,-0.0126390890005429,-0.0297617663359139,0.00428689819320405,0.00397716029709505,-0.0294324463928525,-0.0225787478252779,-0.00935007535553778,0.00178157001672608
"339",-0.00258070484383122,0.00759017276450247,0.00451781769923776,0.0102930540542312,0.00897780571984685,0.00645064661958905,-0.000435233159130521,0.00721911871529235,0.0165462363085529,0.016260283314486
"340",-0.00186815434114684,-0.00599017796499735,-0.0157417474699718,-0.00816399931363077,0.00368912254979703,0.00112484566505189,-0.00711293535248647,-0.00663002781526667,0.00206327377494908,0.015499896788278
"341",0.0112308537949526,0.0114133946489452,0.00380805106175108,0.0128571488475051,-0.00151301782228819,-0.0016852529093877,0.0213451076311622,0.00270573603671109,-0.00491878299974347,-0.0169866569386756
"342",0.000142569404138593,-0.00496527533391056,0.000758397888153572,0.00476857951348575,-0.0109353581966789,-0.00832577794045297,0.0052963345334136,-0.00845447301910596,-0.0183929076535903,0.00550965867879594
"343",0.00206400550283781,-0.00217748991740174,0.00909816692300236,0.00240604071030415,0.000438022894851287,-0.000340563013861317,0.00669217053493787,0.00598660622727598,-0.00222510835256018,-0.0161893475568939
"344",0.0125033038173354,0.0136387581871955,0.019533980035864,0.0212724913087126,0.00908134690825491,0.00556119108618147,0.0124472361940631,0.0126241604200521,0.0211267965185493,0.0113924318653231
"345",0.000912195240340807,0.0123791205718291,0.00368460014610106,0.0127329088304733,-0.00412044137127965,-0.00169227422050444,-0.00656655551638541,0.001958744077178,0.0241379080459769,0.0145181541236565
"346",0.0027334850492462,-0.00301257102689911,-0.00146837588770199,0.000193089220567488,0.00130658804922446,0.00226153707313492,0.00759432144868244,-0.0120864702212312,0.00325478121784029,0.00148039177348736
"347",-0.00810872493699599,-0.00684326105536381,-0.00882381494989548,-0.0173403129920561,0.00521982970443857,0.00304472412878232,-0.0206563019498629,-0.00791642072413823,0.0168923035786139,0.0137964968803499
"348",-0.016914848944697,-0.00912740535193191,-0.0178039233135217,-0.0101679849441251,0.000215783064100528,-0.00236169508078332,-0.0216615101850239,-0.0126952375511012,0.0116611328567406,0.0291615105691487
"349",0.000143421875753225,0.0105662044670232,0.0143503267899385,0.00291618162984908,-0.0117881803905207,-0.0065382654031243,-0.00670059300462389,0.0121234918106492,-0.0106567639262372,-0.0144037392189068
"350",-0.0134043466095929,-0.0119750396416537,-0.0081901881255918,-0.0174452912013764,0.00437749086847572,0.00442478170642224,-0.00645294425444465,-0.0098002567438279,0.00274785658118737,0.00191664407877123
"351",0.00741102905226332,-0.00388923012986098,0.00300243721964488,-0.00161414841801255,-0.00675587798904986,-0.00485723352485357,0.0143175441945003,-0.00751483052741819,-0.0204976645676532,-0.0160210091301101
"352",0.00461580705736275,0.00381365446559223,-0.0112273482471116,0.0134726621270138,-0.00888655092382007,-0.00749237301352046,0.00407474489217274,0.00757173080118823,-0.00246197401004944,0.00631828367677323
"353",0.00502466343160823,-0.00597012896001248,0.0113548329104853,0.0021932873199173,-0.00719489968294784,-0.00468974526054888,0.0104347539032257,-0.00494894936044732,-0.0295041174501247,-0.0272880294777116
"354",0.00250004800066317,0.00200208386185419,0.0134734371304444,0.0034492259470158,0.00657735714098573,0.00333297598672155,-0.00401620479446163,0.00202668219493995,0.0108657378137615,0.00670297976193712
"355",-0.0103312705207066,-0.0148942250438084,0.0022155323035995,-0.0118972589006777,0.00385830686207744,0.00594244838493885,-0.0139688245575832,-0.00845606107566987,0.00583192701538926,0.0133169815653049
"356",-0.00583150142709166,-0.00295030375198546,-0.000736848305582849,-0.0180598672693459,0.00719800460826736,0.00525586582992554,0.000729745629764578,-0.0142753371488895,-0.0122783311991624,-0.023606741866913
"357",-0.000506916095227683,-0.00989345131252106,0.0117993879301626,-0.00871942977938767,-0.00890632448803308,-0.00363697272623809,0.00554624900498468,0.00921574779590206,-0.00264727219085892,-0.0149551263085738
"358",0.0199972440145992,0.0193311974814387,0.0080176690744489,0.0318167539879337,-0.00599023861740622,-0.00524760744759589,0.0251088764717735,0.00913152031209297,-0.0023081938301629,0.0379554310072467
"359",-0.0318936703750909,-0.0281265831677109,-0.0354306334481762,-0.0362303416298275,0.0129464051276929,0.00871614780441443,-0.0396429652400664,-0.023268833203281,0.0301908743848771,0.0255972879346751
"360",0.00242110407008589,-0.00103678910035232,0.00149919667326714,-0.00255702560647619,0,-0.00716279480465831,-0.023146459342973,-0.0138019950188428,-0.0120143726030624,0.0102211742407385
"361",-0.00497708954951881,-0.0136831297723301,-0.0217062658025592,-0.0230705077771063,-0.00650080470056469,-0.00595444082064356,0.00392417226802677,-0.0279905751162335,-0.0277303677174762,-0.00400007566573857
"362",-0.0147124943588905,-0.0154996561237104,-0.0145372347765824,-0.0149635932726708,-0.00232907953453321,0.00103698501317373,-0.0205954811368967,-0.00394509718179681,0.017182863219771,0.0368531702795376
"363",0.0038076922212682,-0.000874241415392496,-0.00232906154917489,0.00583161343547212,-0.0100041363377068,-0.00874600596359998,0.00613995523585187,-0.0128711167336001,-0.0163180768668609,-0.000227787839221172
"364",0.0126439829890479,0.00787878365522676,0.0101165083611312,0.0108082340738569,-0.00213365857386905,-0.00232200952549866,0.0208996681774209,0.00902712645860992,0.00268696267960178,-0.00638108513231939
"365",0.000587817995276074,0.00550092647301526,0.00924517614482756,0.00339914327566926,0.000225719457783491,0.00011628566338473,0.0143457817837016,0.0069582287762513,0.0137481064022347,-0.000917259715971785
"366",-0.00484499494108648,0.0012473539233786,0.00687002772180811,0.004234063358314,0.00202540399818107,0.00337404074323033,-0.0294639421882777,0.00592292736706757,0.0027582805939943,0.0101008964033154
"367",-0.00973621360897714,-0.0107362890590078,-0.0106137209988637,-0.00484900165369406,0.00841937273879223,0.00545035812006356,-0.014875540455104,-0.0107951224702459,0.0118051461318052,0.0136363564003168
"368",0.00126605254689593,-0.00164708260652724,-0.00306509293330259,0.00155386126818668,-0.00590027910761159,-0.00576624993922858,0.0206470049094201,-0.00297607663388588,0.00158585185303406,-0.0233182687419895
"369",-0.0162318738245886,-0.0198000405545667,-0.0330518426047427,-0.0326449420222619,0.00582340374408452,0.00463933783566239,-0.0247582027116291,-0.0107121542683088,0.00599410780353082,0.00688701191158803
"370",-0.000987966545401231,-0.0037210041200606,0.00715410106663428,0.00291527238845246,0.00211663869251288,-0.000460992172904517,-0.0207427840733845,-0.0207612264464411,-0.0209106358935571,0.00706784901461277
"371",-0.00197796539858042,-0.00377541853317043,-0.00789228111496521,-0.00443297162141409,0.0066652404481724,0.00531330870924585,0.000473860696870165,-0.0022866603377284,0.00436335994320181,0.000226438523680317
"372",0.00472579575528265,0.0134181607292101,0.0151875664578527,0.0200241362875024,0.000441980106322015,-0.000116233646972441,0.0176525160989316,0.0177083408968977,-0.000571658847928758,-0.00384796818793998
"373",-0.0271600708997232,-0.0245604227631595,-0.0251966634692354,-0.034310549460141,0.00672970978020793,0.00563213972865739,-0.0357588910249208,-0.0227228009415239,0.0364905407570473,0.0331744203459301
"374",-0.00545880790453213,0.00466275090232049,0.00565388658704746,0.00966900129928239,0.0117265818253598,0.00491339621463904,-0.00780718138147207,-0.00691238024990404,0.00949122602923258,0.00263902291314744
"375",0.00352844535824359,0.00268134775606277,0.00160667547620763,0.0075728474254606,0.000216103949540303,0.000682012149010758,-0.00327900233775269,-0.0101242841182188,-0.000765267292388017,-0.0177670229074153
"376",0.0031254150494644,-0.00874297843131866,0.0040097357658313,-0.0178311591764355,-0.00236930166058535,-0.00271341680027215,0.00575666747909986,-0.0100149385494493,0.0137855795670552,0.0176417854465454
"377",-0.0171366053934826,-0.0153574568132856,-0.0215653831264279,-0.0285067418969485,0.0052294058626019,0.00240120854446624,-0.0207684201180174,-0.0079636807646134,0.00550392810257172,0.0190915051542797
"378",0.00103056332151241,0.00779861350377642,0.00326514509197073,-0.00285762647823717,-0.00216803032313317,0.000342551117810563,-0.00801644438086335,-0.00282072284157864,-0.0119137063843235,-0.000430672741844051
"379",-0.0102129881570902,-0.0119210694509649,0,-0.00356216020008893,0.00456198320641565,0.00467364337699538,-0.0205383403951658,-0.000217683188597384,-0.00901580510570943,-0.013571687391414
"380",0.0177569287154768,0.00910150828758272,-0.00406816674301513,0.0122795736137693,0.00648788033508385,0.00249676966065038,0.0723612897245027,-0.00217604168830665,-0.00405570522671139,-0.0362524577358925
"381",-0.0192548508598467,-0.00985845931076734,-0.0163399534131995,-0.0201919820434368,0.0044042837583238,0.00475432642475515,-0.0735695695479364,-0.00719723112665738,0.00704379257050647,-0.000679765429519197
"382",0.00408696796583485,0.00646107647417882,0.00913604548925417,0.0181007629802203,-0.000107358923278067,0.000338159403751037,0.0181659478003791,0.00395391639049003,0.0221857814207651,0.0272107961405996
"383",-0.0116520826722747,-0.0181013367537142,-0.0131687754605394,-0.00669595684399071,-0.0142259811370272,-0.00934737104583483,0.000340255182767368,-0.0205687226562405,0.0174276169937733,0.0139072576091852
"384",-0.009044222752426,-0.00321534750206998,0.00667260657963009,-0.00123984400322441,0.00878898848046417,0.00534328106286175,-0.0348223632361876,-0.00379792257377121,0.00788146246820243,0.000435523166912199
"385",-0.0140969052911251,-0.0148387376178717,-0.0165701926879738,-0.0166798442948501,-0.000322484003253631,0.00361789636804133,-0.00950390075786112,-0.0222026428657347,0.00271081210673296,-0.0317736170793276
"386",0.0245472641234239,0.0128791333448321,0.025273537219308,0.0288760418543093,-0.0180761807593485,-0.00912630578206208,0.070184921177403,0.0155964541340976,-0.0179889366328155,-0.015284340931413
"387",0.0100032424285166,0.0223062339032079,-0.00493007637350207,0.00467740704386443,-0.00515090729080658,-0.0047765225443237,0.0161046618137299,0.0219058089178112,-0.00232953192864194,-0.0235107378302527
"388",0.0062301791513224,0.00980274327051434,-0.00412863539291763,-0.0086245234447262,-0.00374530043756716,-0.00342729688155075,0.000326895651196812,0.00773499292244129,-0.000530704727969455,-0.0170640232062798
"389",0.000555602650132547,0.00584570118755967,0,0.0123953174353453,0.00387113356098578,0.00229296533986556,0.00294043120301368,0.0164471913093296,0.0100881917826949,0.0121285500252375
"390",0.0113444717088964,-0.00010416882207076,0.0132673240537253,0.000608215169020765,-0.00495698308986958,-0.00343168554766515,0.031758956461087,0.00539390891588676,-0.0216569063817208,-0.0218516034181685
"391",0.00541308044894606,0.0035291308127765,0.00654614703337808,0.0014440080293745,-0.00199185187582551,-0.0016064257516446,0.0213099184780294,0.0313304269854897,-0.0267569100957857,-0.0225799169704837
"392",-0.0207539222231441,-0.0212015989251964,-0.000812912871918647,-0.0369583531770727,0.00975899190832963,0.0086223111282524,-0.061514612970518,-0.00728249617207444,0.00839132162967871,0.000737439518115224
"393",-0.000239226546505322,0.00612827005524896,-0.0113914432196633,0.00685547477954929,-0.00999395888227483,-0.00581342336518476,0.0151515686414065,-0.0253613140873827,0.00394174961257554,-0.0125246920014604
"394",-0.0146636478184291,-0.0149129196484419,-0.0115225290458678,-0.0169051803573517,0.010094846361737,0.00573262589743373,-0.0212525550043362,-0.01096762757253,0.000436263487048283,0.00497402307860817
"395",0.0213526062335463,0.0110875368600938,0.00582837228450406,0.0554093630688424,-0.00406294780344074,-0.00285032230288906,0.0500582812305685,0.00217423237812708,-0.0124278530765991,-0.0113834159100783
"396",0.017817604308429,0.00991126217869231,0.00910609586463718,-0.0104094139742621,0.000991788811586236,0.00194453763091862,-0.00489344666221658,0.0197439256027891,-0.0118114477011346,0.0197747231077408
"397",-0.0132265967106729,-0.0110667414340564,-0.0155865551292548,-0.0224103921468032,0.0099154738084446,0.00798630875330231,-0.0117388340699155,-0.00531931043827449,0.00625564140713708,-0.00834558517007378
"398",-0.00528294556007392,-0.0130912920175436,-0.0141668964883657,-0.00678379215505653,0.00221168810835981,0.000499870033491501,0.00240790318608597,-0.00342241857290793,-0.00566165617980341,-0.0111386394825681
"399",-0.00927392374367209,-0.00363738855405171,-0.025358896777375,-0.0306163819642299,-0.00229423751633739,-0.000680677958422859,-0.0140914189806951,-0.0223224072682821,-0.0159651780730155,-0.0330412197272842
"400",0.0269622066986863,0.0300623017804762,0.0225497678284565,0.0128762119076171,-0.00744538134200778,-0.00511263236182546,0.0427155581139227,0.0208564385968686,-0.0233718745560686,-0.00698947251736459
"401",0.00444083022089181,0.00145940412514123,-0.00593723137353508,0.0199089981193943,-0.00408154446927711,0.000342147662914405,-0.00467287468555388,0.00559157877414496,0.00650554120572644,-0.0106882484373897
"402",-0.0148917213399747,-0.0185264790108302,-0.0221842795380595,-0.0343370064215143,0.0162822858187175,0.0093613958839005,-0.0242567726250514,-0.0248079629295906,-0.00634814180918908,0.00553359520466379
"403",0.0185812823596383,0.00042438831899716,0.014833917411067,0.00243591150588807,0.00272490486599031,-0.000452373418758145,0.0323978660421715,0.00197372410256746,-0.0192821010236776,-0.0280398631922217
"404",0.0103576783187704,-0.00190766920883678,0.00601901864658161,-0.0104474923013772,-0.0095653516251718,-0.00486625659352213,0.0245453231651027,0.00656633252370664,-0.0390856686012081,-0.00107836893611957
"405",-0.0104045379286555,-0.00488566245456112,-0.00683768511669636,-0.00834757076741366,0.00932857931260567,0.00693579589712567,-0.022137721984121,-0.00478405222738409,-0.00751879727050897,-0.00863694178083629
"406",-0.00603014263486812,-0.0175026428880108,-0.0172114074098775,-0.000247616070586654,-0.00347924702567226,-0.00214477893318876,-0.0161265836961962,-0.0190080454938174,0.0129160586034298,0.0334875668411299
"407",0.0075443577214267,-0.00695187274977271,-0.00612946058170472,0.0131252885364186,0.00643680038087036,0.00305454329118349,0.0165486938781636,-0.0144764183357673,-0.0270966166526879,-0.00869334665424149
"408",0.00486349924375706,-0.00700063308171139,-0.00704874966022784,-0.0156439029518063,0.00867363406307575,0.00372331654653246,-0.00155026991268004,-0.00338998581073546,-0.0216761316112446,-0.0135530788405448
"409",-0.0136743651509919,-0.00638938058928429,0.00887314830507457,-0.016885907937036,0.00397634672918601,0.00247323068331373,-0.0209627781349175,-0.00680294599674813,0.0150715708516644,0.00565732592459312
"410",-0.0109041585400537,-0.0121949744562655,-0.0158311411676602,-0.00833589863150708,-0.00385434758546832,-0.00145808697196048,-0.0206184694768672,-0.022830911349251,0.0206852403292421,0.0155371930081818
"411",0.0046456540547386,0.00224485358181403,0.0107240905599848,0.0254713512586842,0.00279490566847285,0.00291998767330992,0.00242892526993077,0.0163553052918237,-0.00460029839612097,0.00791332262534139
"412",0.00172451399668572,0.00515082356113594,0.00618878012850099,-0.00148995438297961,-0.00182141749504094,-0.00212765064718912,-0.0137318811290084,-0.0114945132943785,0.0279790788903094,0.0429208050077479
"413",0.0144754815028982,0.00713013501557325,-0.00702985182691929,-0.000746803915695926,-0.000644270779306511,-0.00291722022651242,0.0229321612298448,0.0090700419653349,-0.0148238269201523,-0.0338770128588113
"414",-0.0202850342443994,-0.0163716634029967,-0.00884929794196343,-0.0206620575629712,0.00999124352309111,0.00663876619831716,-0.0220981071301368,0.00230473961868682,-0.00185004928835575,-0.00571443886543999
"415",0.00291280531299809,0.00382382626462618,0.00535694647780538,0.00177977035499888,0.000851315375291151,0.00033581918100456,0.00769625846262612,-0.00436896718114477,0.00370694427282814,0.000522586882356402
"416",0.0097335185499654,0.0109791746544148,0.00444083723943867,0.0213140165558947,0.00170059254423438,0.00145218179033324,0.00893775709393196,0.00808342302194798,0.00160036926257412,0.00939941240979691
"417",0.0121283278463378,0.0141845724471144,0.0079569991989259,0.00695673129236529,0.000105877234568785,-0.00145007601634783,0.0331769327216458,0.0119127074527881,0.0100786503186008,-0.0196584834087645
"418",-0.0107535466379791,-0.00611914046883755,0.000877488672929472,-0.0118435055404527,-0.00445585587555386,-0.00122864783664056,-0.0112234752467776,0.00271665536991827,-0.00571916524701888,-0.00369406808285622
"419",-0.00621160583876113,-0.0127528497788023,-0.0131464395913908,-0.0302119210926047,0.00930477574423416,0.0054434927836049,0.0122971837419723,-0.00541898375988015,-0.0307184191741331,-0.0259532462648115
"420",-0.000859765781231481,-0.00467690271026078,0.00444083723943867,-0.0164778497819016,0.00423789898792193,0.00245629339592401,0.0137046130228049,-0.00726420998991073,-0.00391411630987804,-0.00570970809837212
"421",-0.0301059875127838,-0.0449766273421935,-0.0318305929064672,-0.0460732670500286,0.00802023572047061,0.00501161212730672,-0.0311872180350191,-0.0420764419771621,-0.00633793898260793,-0.0142191914588167
"422",0.0031442354448632,-0.00562315817243786,0,0.014270009993067,-0.000523369793648754,-0.00221664528858279,0.00634304776488159,0.00501309214160872,0.00752652133596787,-0.00998620532375682
"423",0.0206560884282787,0.0172008825832166,0.0246576310382751,0.0124460139694795,0.00418886861647239,0.000110885666798177,0.0431771777822469,0.0261284571030778,-0.00151939725806294,-0.00224151519185878
"424",-0.0296876410782867,-0.0277971192717003,-0.0276293663373014,-0.0561200332085667,0.00990818954739514,0.00455331570537765,-0.0438068010335202,-0.0199073431015574,-0.0300532966008965,-0.0365066424621719
"425",0.00405787011146108,0.00428872942971847,0.0128323703816309,0.0161383169800058,-0.00619597552020679,-0.00254194567310118,0.00537123342963408,0.0243269671110884,-0.0296770435266582,0.00145725716199618
"426",0.0144680233760981,0.00142338148894505,-0.00542977565125347,-0.0147672495141199,-0.000520137449865565,-0.00177337795819965,0.0114706460508218,-0.00807024010396307,-0.0153597276292141,-0.00844003600158705
"427",0.00462113472377679,0.0234543697946199,0.0063695334162186,0.0333708586139994,-0.0128920373412226,-0.00499682020134384,0.0105640017535407,0.0167364218239567,0.0337985896606847,0.00675078805886775
"428",-0.0475848203942226,-0.0467593312533753,-0.0280290632558463,-0.0785441558822995,0.0324409503723111,0.0191930223361763,-0.0614911781634634,-0.0477824947542697,0.026604830181145,-0.0393584528508193
"429",0.0167371015520763,-0.0118991307965071,-0.00930247357594216,0.0086131444139439,-0.000204218085122498,-0.0028468018837563,0.0307945468197177,-0.0177671241212914,-0.00992775941020507,-0.020333922337049
"430",-0.0449628722150951,-0.0459568995708661,-0.035680664758161,-0.0709658021308874,0.00500094264847917,0.00900274590190575,-0.0465599294224486,-0.0381325454457248,0.11290529869898,0.0300495994542949
"431",0.0296713224254774,0.0569291622921919,0.0447907663797411,0.0843106421454241,-0.0146208960728207,-0.0117515611887198,0.0845002940384527,0.0200763663933543,-0.0311256263880836,0.0018046140202741
"432",0.0397140871234507,0.0714108415443078,0.0540542568663878,0.124525084458892,-0.0317364267568371,-0.0178385034174465,0.0327339562995848,0.0652989271150723,0.0384057957099349,0.0330228692629901
"433",-0.0226395683224588,-0.0204729344068474,-0.0344829616581471,-0.0652458500917913,-0.000106155125931373,-0.00212954424739209,-0.0880951430125682,-0.0179792483670932,0.0372179214741364,0.0345829335306627
"434",-0.0227515430511512,-0.0234552869030249,-0.00915776543959201,-0.0311454849646861,-0.00383183110046326,0,0.00636379160417633,-0.0158998080893874,-0.00964341780668332,-0.00983125370641769
"435",0.00320527141008298,-0.0019027273124772,0.0138633000910231,0.0114811275784215,0.00438050496806031,0.00258458165406439,-0.00739000328331385,-0.00612064515083111,-0.0182291779891304,-0.00822696864585204
"436",0.0156394418493786,0.0243030941927633,0.0173200594729372,0.0513618202767543,-0.00202088631351416,-0.00302579114101509,0.0185308768956625,0.0187197375565189,-0.00299852384959665,0.0174484640515546
"437",0.000496636726029731,-0.0093045575148093,-0.00537655465979003,-0.0340080871140672,0.00724780405371184,-0.000674468308489939,0.0207925805946605,0.00580240269627108,0.00219782540883151,-0.0118076703580804
"438",-0.0783614064740071,-0.103545610456054,-0.0774774377757225,-0.116792296379982,0.0291003652931663,0.0139463632252481,-0.0598344922335913,-0.0973555490220709,0.0338181098086114,-0.0620198269049511
"439",0.0413896891885062,0.0440025932392998,0.0410157898931347,0.0809868257571509,-0.0243697804467896,-0.0131995454376148,0.0485781856703116,0.0162449283182604,-0.0502400357262476,0.0279040396033075
"440",0.000603431226825712,-0.0012549039672608,-0.012195225838988,0.0119989779034817,0.0125801280638027,0.00704929756444761,-0.0153347513177419,0.00943414444230495,0.0105795345009991,-0.0233106248146986
"441",-0.0362742150570512,-0.0419491843303595,-0.042734953546995,-0.0876229280186489,0.00803923662701234,0.00560093709329901,-0.0662299230647353,-0.0501041215787444,-0.0423403391608662,-0.0552870733393158
"442",-0.013500170888456,0.00209779020492284,-0.0198412566138197,-0.0263074410885342,0.00880409372558999,0.00378678171761826,-0.0533705705148634,-0.0213173477157439,0.00315794963784888,-0.023345023034933
"443",-0.0509335360088863,-0.058084873512945,-0.0323886664484032,-0.0751951604800709,0.0181722618067408,0.00809983605722375,-0.0183605250165393,-0.0823790818693318,0.0204625630445605,-0.0425672076916122
"444",-0.0447860929286437,-0.0500000731876666,-0.0366107034530171,-0.0777896710539274,-0.0030252225148909,-0.000769960164404893,-0.0844511904582392,-0.001826138199711,0.0354769581807897,0.0123118879564208
"445",-0.0251925978017469,-0.0102341143502516,-0.0369164653807771,0,-0.014362220545762,-0.0127783340471617,-0.0167151084771379,-0.0423780788829878,0.0246361988530834,0.014527083835969
"446",-0.0698389573512856,-0.0747412186942116,-0.0462232272372948,-0.073663989320263,-0.00841429255722981,-0.0100414185369551,-0.071562977533294,-0.0799106929849241,0.00536797149111989,-0.0466200320130208
"447",-0.0242556946137834,-0.0249043592518915,-0.0437351742147506,0.0115368008871644,-0.00703730068428776,-0.011723439996784,0.0795657473149818,-0.0311418098450797,-0.074304792562741,-0.0443590389076348
"448",0.145197732346766,0.137524774725515,0.158220049558436,0.227698446195007,-0.012819029863942,-0.00684277107973541,0.074748617265141,0.107143081748968,-0.0147801368086982,0.0555555194676047
"449",-0.0148000952855143,-0.018422792685358,-0.00533632816919272,-0.0497675591118867,-0.0064405851438063,-0.00470819714297233,-0.0648741927635226,0.0438709627228235,0.00256127582781485,-0.0183518618979334
"450",-0.0984478872247684,-0.105571683876009,-0.104077164913132,-0.161662192913883,0.00956385110213365,0.00819183742345975,-0.141666651800415,-0.0908531636396415,0.0135036622933209,-0.0455026021484503
"451",0.0416572698355069,0.0498358069609481,0.0610777823579713,0.0491463009638773,-0.00515731543467546,0.000228893915418027,0.0628639998588265,0.047246928907658,-0.0482534761314001,-0.0188469788539656
"452",-0.00597204498315018,-0.0162397112971843,-0.0135438985971369,-0.0313614985660879,-0.00687737562584234,0.00629293975048872,-0.0102764984269611,-0.0327815538009583,-0.0262328411371821,0.0112994087772322
"453",0.0600798490158407,0.0520634605726538,0.078947104108916,0.0700817106203804,0.00798964712447092,0.00102322036751157,0.00946014659426675,0.0620804900339498,0.0167076935203692,0.0201117479402557
"454",-0.0298553391095193,-0.0585395150052697,-0.0360549633603064,-0.0796630898511226,0.00528459096038003,0.0105633974240107,-0.0345142325024468,-0.0423380226274573,-0.0314649808917197,-0.0357795082209367
"455",-0.0544542741607011,-0.0762821727153007,-0.0605061097692504,-0.105284984649677,0.0202902720743121,0.00764343056252259,-0.073390130072325,-0.0514680790064955,-0.0568196771908416,-0.0473305935845669
"456",0.0115840176859305,0.018390024720764,0.0339580451129045,0.0279070369975749,0.00741919699102378,0.00133902710317813,-0.0155853568488339,-0.0285219746789565,-0.0147817182370898,0.00397460927152582
"457",-0.0507142206187731,-0.0494035228559396,-0.0600226604224522,-0.10316762595156,-0.0106376465205411,-0.00423369159962594,-0.0641057654766138,-0.0748298527207426,0.022080636317604,-0.0399841171555951
"458",-0.0355008936122312,-0.0580645787019431,-0.0602411813573567,-0.0262358983086028,0.000723842671334296,-0.000559697476548937,-0.0521350662971245,-0.0170280197192976,-0.000415441080396484,-0.00742275787031688
"459",0.116855442870684,0.129756344945488,0.121795029265195,0.209326404702385,-0.0145658323937473,-0.00805906614240925,0.16325336733421,0.0362206249324153,0.0223053615960098,0.0274200670797233
"460",-0.0072530238366737,0.0148199019911786,-0.022857192870795,-0.0317050240210727,-0.00503227738998269,0.00146685217153641,-0.0397386835719666,0.0136780030800543,0.00284590048995925,0.059037684233568
"461",0.0345939786823455,0.0288749474849697,0.0538010882657642,0.13495604675344,-0.00906090035008733,-0.00766169956165097,0.0484549605510589,0.0468512987598091,-0.017432445945946,-0.0412371829495353
"462",0.00550362467139909,0.0125804886927852,-0.00110988216421792,-0.00857748700177363,-0.0129726912342244,-0.00204353321365069,0.0629526693993792,0.0204081478810851,-0.0188420164879936,0.0111509323669647
"463",0.00289171770462571,-0.00382290684292108,0.00666655769421842,-0.00904427751586756,0.00270451643308944,0.00159838790655509,-0.0364278717371116,0.0245614996523509,-0.00336414372661309,-0.0110279603272104
"464",0.0339821855694262,0.0697155290151585,0.0551877219015868,0.0912697513390806,0.0187681515730052,0.0119717043812242,0.0556098441367348,0.0352737580864686,0.0616034475837819,0.0454003257497158
"465",-0.042027655355218,-0.0594919043279867,-0.0209205195797366,-0.12727260225598,0.0118586863483465,0.00529409623446009,-0.0965801906426051,-0.0370491467601426,-0.0355060929184117,-0.0259048539988933
"466",-0.0554112648199867,-0.0632547519414924,-0.0865383446173636,-0.050416866206113,-0.00722076700435215,-0.00302510694747138,-0.0452690646729317,-0.0398483500573027,-0.00796706011124759,-0.0438013163797875
"467",0.0330176159397382,0.0563285731220824,0.0584795746067168,0.0811759961838443,-0.00653421868010173,-0.00359744516784133,0.0592023491856679,0.0296949160249347,0.00387702847027116,0.00122699958366002
"468",-0.0131043069526336,-0.0215227337317717,0.00883967803428454,0.00933440741949076,0.00487991738568549,0.00101606750390459,-0.0857363682871138,-0.0535088668463697,0.0148965793103448,0.00653592119552315
"469",-0.0308757207054389,-0.0252792277379935,-0.0416209230279155,-0.0623241473770969,0.00295656338472838,0.00371860041433925,-0.0127247797493318,-0.0326726541377507,-0.0207936797827213,-0.0190745666179768
"470",-0.0440011898211417,-0.0565845788383202,-0.0274287421471091,-0.0741851059680003,0.00642065721734086,0.00617531709392494,-0.0736900530970118,-0.0288422886190112,-0.0284525040200208,-0.0293754072624588
"471",0.0623395085318368,0.0828275950225159,0.068155269169891,0.138489850314846,-0.0239516762645893,-0.00725321910867283,0.110708229457389,0.044157722414307,0.0307143142857143,0.0187553871036426
"472",-0.0499064178101235,-0.0524234748979634,-0.0539053251836887,-0.0960129816234701,0.0198242790378005,0.0098917006770125,-0.0985839058187041,-0.0550149569772006,0.0159390293571995,-0.00627609242624128
"473",-0.0132763220224886,-0.032706875247617,-0.00232558990830822,-0.0166512138976598,0.00441329883756314,0.00422996766480921,-0.0078550504576691,-0.0213863993173454,-0.0088676804010499,-0.0227369028419511
"474",0.0188369360605409,0.0143883900657971,0,-0.0146456180382868,0.0128677311700669,0.00775890596911455,-0.0401949764507754,-0.0129499851238185,-0.00192704743490579,-0.0150796573222827
"475",-0.0640789426184306,-0.0606380766249911,-0.0641027640217685,-0.0863912897266207,0.0256140989253113,0.0107778423872322,-0.120558376285,-0.0873311466723421,-0.00344780020830782,-0.0113736460813515
"476",-0.0742332575120096,-0.0683278371020931,-0.0286425507123564,-0.0716825088598804,0.0516619712046136,0.0201317265965206,-0.0873018639228385,-0.0336921791110484,0.016468239234203,-0.050884855047417
"477",0.0539425094417376,0.0571313521477923,0.0615383098893156,0.144030350549349,-0.0144596086303003,-0.00917320490438767,0.082609008565327,0.0418406441548014,0.0735194175705685,0.0172494312916369
"478",0.0692913901329324,0.0770407259505146,0.0471016369669053,0.06079468372803,-0.0156435121544644,-0.00936699360873539,0.144578188882891,0.0441767092283893,0.0261256316074987,0.0687441540990277
"479",0.00740914148088723,0.0202850149180385,-0.00461383718925945,-0.0189531213551635,0.0294150307743162,0.017170763102166,0.0271131367046289,0.020940113368118,-0.000494388802650403,-0.0334477063449429
"480",0.0386409421501512,0.0177883948349757,0.0185402269866948,0.0763573470976295,0.00134252146638825,0.00608996292987785,0.045652447042692,0.0397658580076123,-0.00605918117747561,0.0319432230558587
"481",0.0125886945934564,0.00342718915434892,-0.0147895207106529,-0.0192309687276792,0.0123529473873265,0.00201689556376028,-0.00861300958211364,0.0362318086785434,-0.000870850990452365,-0.0434221329352545
"482",-0.0885780296579917,-0.0877732942633797,-0.0577368686040384,-0.0962962868118226,0.0382949084254187,0.0135358618188552,-0.206111689351636,-0.0784771274728431,-0.0580251041719612,-0.0310112387636797
"483",0.0384848141377605,0.0490450605743009,0.050245035940212,0.0631625615563265,0.00383947936841422,0.00524595793603733,0.137735930385694,0.0408939316547603,0.017184335302463,0.000463807880641598
"484",0.0240413406304854,0.00749459841093225,0.00933499704839735,0.00816367917750171,0.00282256941651982,0.0015652633629033,0.0454396774480499,-0.0064805063469735,-0.0100064591295564,-0.0115902577741106
"485",-0.0231333659476316,-0.0262128164843534,-0.0393061261241021,-0.0427351675050608,0.0197042479283107,0.00625152626808667,-0.016497397270961,-0.0342438197670699,-0.00892622735626158,-0.052532722436711
"486",0.0308321145295809,0.015278126759841,0.0156435317965196,0.0592108699575564,-0.0162062652294602,-0.0105616752138862,0.0964516194263618,0.00253284399542508,-0.0129801721854305,-0.0247524516760373
"487",0.0349141626528939,0.0458616494271007,0.0450239085583943,0.0638859968294161,-0.00217263364743192,-0.00376736443234771,0.0941447051856283,0.0484211230425975,0.0225442843214285,0.0461928228227908
"488",-0.0164835166378312,-0.00548145780909037,-0.00680284926262409,-0.013761381373292,0.0197751112756526,0.00850933954068678,-0.0717929453658296,-0.000803433208772519,0.00170610242937408,-0.0218341123036047
"489",0.0068155644700274,0.0285913424588287,0.0216891662498477,0.0596195024432267,-0.00240231519320644,-0.000937741151985749,0.0663382816060714,0.0478292514823961,0.0448054226436416,0.0302580101527612
"490",-0.0240811657343912,-0.000669837823792152,-0.00335159721632461,-0.0255384920651915,0.00196203058351974,0.00604700359310617,-0.144254340756472,-0.00460234832389383,0.0112852915360502,0.0317765472120874
"491",0.0119394597721407,0.00502676923333922,0.0224213384009773,0.0139230783678752,0,0.00279860156527323,0.0946030616987708,0.00346805281583551,0.00198383132092173,0.0219319417556862
"492",-0.0139339515555288,-0.00200089782537349,-0.00548231202183491,-0.0133283749012244,0.0113907512660145,0.00217018195499419,-0.0284223327345389,0.0145929688930451,0.0221507244685244,-0.0282931297013179
"493",0.0470655240948976,0.0648180932727804,0.0507170765587521,0.0798201248114623,0.0247247753348434,0.0158810414482828,0.121791095135272,0.0264948865507211,0.0225181724580672,0.0143198584309669
"494",-0.0096866223188361,-0.00972705195447299,-0.00209896071555626,-0.0174372425870895,0.0271344651554184,0.00680154384215559,0.0252792580410466,-0.00921813799145765,0.0114847384736532,-0.0136472101417828
"495",-0.0186831692398535,-0.0323193797957069,-0.0347004776186026,-0.0219909383607423,0.0209827172006971,0.00675518851754031,-0.0788992488363667,0.00446553420223506,-0.0182605290881425,-0.015267213431192
"496",-0.0043017957093987,-0.021610933434199,-0.00435715070259834,0.00355032317496584,0.0010650653553117,-0.00330476193629659,0.0495912179124531,-0.00156732464611442,-0.0147848569887377,-0.00678285373721177
"497",-0.0128133705375975,-0.000576063938044769,-0.00218839077867405,-0.0373428248206685,-0.00768871870728738,-0.00261271013901043,-0.0209395191737293,-0.0332709756759678,0.0100448024946678,-0.0282925977976181
"498",-0.0103374320363466,-0.00576477054041391,-0.0171363780834707,-0.00828142206825622,-0.00131920595129442,-0.000503742280340447,-0.00759272884242845,0.022814758170411,-0.0099449078593925,0.00401600906206068
"499",0.00580277875870228,0.0133013567625655,0.0123735264415281,0.00709800599220234,-0.0021461301828879,-0.00100849089347121,0.00765081943985768,-0.00189029629703064,0.0100448024946678,-0.0154999422095188
"500",0.00576987124169337,0.00807828959965962,0.0188889991519015,-0.00331654255531411,0.00330891673902634,0.00534874538572461,0.0132173908266688,-0.00378732075196853,0.0256410139664631,0.0157439728792961
"501",-0.00286821815909899,0.000333688716982472,0.00763336961302619,-0.00166420856781002,-0.00119946348341327,0.00220582226089472,-0.0563420469884768,0.0112015040428302,0.00876168244770281,0.0110000038080995
"502",0.0237026429906173,0.028371260668163,0.0281384680100631,0.0266665798747225,0.0095236402851393,0.00140678692114404,0.0452940609293955,0.0113036081756854,-0.00521130295799199,0.00593463684071205
"503",0.0142743306334083,0.0107109315664768,0.00842097678856013,0.0133930591584175,-0.0209187105269434,-0.0110403101491199,0.0475519320091706,0.0089417976746875,0.00721763661891428,0.0417896661742048
"504",0.0301420438654938,0.0105971974697197,0.0052197084709853,0.0476571778360306,-0.0251362753947457,-0.0143104904984849,-0.0273971976728643,0.0347118605047498,-0.00335175693545164,0.0349221404623925
"505",-0.0011834829136359,-0.00953282341030859,-0.0249224444998591,0.012996780845002,-0.0257840264641591,-0.00175100866198741,-0.0196079506217892,-0.0071380908109151,-0.0202945603515751,0.0104879131647666
"506",0.00667748451896255,0.0121911766364733,-0.00958500897038983,0.0226417638325778,-0.0100574484984624,-0.000618437156042484,0.049577578240682,0.0273187336443235,0.00769405749192509,0.0261732517063458
"507",-0.0299560021709716,-0.0117274418778813,-0.00967709258919836,-0.0575645572555606,0.00392113325428189,0.000206469592025416,-0.0338166516334358,-0.0129457741418092,-0.0279572076103797,-0.0510114152463199
"508",0.00408073574899559,0.0128288592182748,0.0141150782402482,-0.00430713179987074,-0.000798989567391106,0.00268274771935739,-0.00444425229188961,0,0.0206646404833837,0.0037070854943253
"509",-0.021419257849012,-0.0345157467355991,-0.0171307549928315,-0.0216278758451942,0.00151070204262282,0.00463093870691211,-0.0460381091495752,-0.0212692980783469,-0.00639357099684534,-0.0115419980752803
"510",-0.0240210173052431,-0.0272216558075102,-0.0119821858531877,-0.0422028342502593,0.0103790678111491,0.00624877143903224,-0.0582038500676512,-0.0315100881933605,-0.0376548626705163,-0.0453058901349086
"511",0.00184053404075391,-0.0188806521965705,-0.018743248956921,0.00293759501993507,0.0010529437440252,0.000712112486840999,0.0301240574750288,-0.0373973281129588,0.00148582215240656,0.0166340748254159
"512",-0.0314541333323711,-0.0474231071146841,-0.0292134512336298,-0.0485353332614654,0.0164887248748955,0.00559559052458836,-0.0518539826999515,-0.0470087229818827,-0.0134767067313318,-0.0139557828393829
"513",0.000354990882136974,0.00649360533073629,0.0127313121313088,0.0114332418117733,0.00163889421160235,-0.000809437400665303,0.0289349509087704,0.00163096426626863,0.00751971415566222,-0.000976072559683128
"514",0.00782004930862024,0.00143373584165674,0.00685749258322121,0.0108695598587198,-0.0154191969654682,-0.0092127199705988,0.0367735555671418,0.00488399960735375,0.0288593112185509,0.00439661793669699
"515",-0.0527861274911735,-0.0776663211707042,-0.043133080226246,-0.0744083209295803,-0.000174413626271352,-0.00153364944641332,-0.108196380926381,-0.0810042145617409,0.0218836660849193,-0.0311282811770387
"516",0.04319218174729,0.0364761653506118,0.0438911610345296,0.0543680991120288,-0.0315896121186571,-0.00890378902901501,0.0995986413544672,0.0599383022351483,-0.00437760308959789,0.00401600906206068
"517",-0.0154669378417212,-0.0243352335811523,-0.0250002771842245,-0.0330545137199784,-0.0192461098635481,-0.00660887449654735,-0.0507601610580918,0.0112262019820739,0.00510992263553356,-0.0129999764309525
"518",0.00435045697077219,-0.00652325704769396,-0.00233073619696078,0.0127622024042979,-0.00783106461350314,0.000208368506275036,0.0317004463462636,-0.0143911220469064,0.0467013112626791,0.0466058108368732
"519",0.00685832541427089,0.0266512433752151,-0.00116844132431437,0.0117012054335544,-0.00872866351231738,-0.00249457747574278,-0.00837990656897025,0.00709187319457971,0.004744131986266,0.00193618162824372
"520",0.0101579500965925,0.0161775683666319,0.0315788867531512,0.0177936042784008,0.0235128147396142,0.00656459290268674,0.0181536803629661,0.00289974871672105,-0.0064080946512004,-0.0270532163348416
"521",0.0338336262323466,0.0373934241901301,0.0181407310453101,0.0506994938112106,-0.0249865991488234,-0.00641834007968534,0.0796186430069112,0.0177616305798252,-0.0108621750688677,0.0238332003545942
"522",-0.0324974133649691,-0.0456815511310791,-0.0378619337583482,-0.0507487969011498,-0.0229980862797431,-0.0130220760438345,-0.0783031998855278,-0.0300324282445924,0.0237932057605399,-0.0121241352363949
"523",-0.0203433796210799,-0.00710580860485432,-0.024305661846818,-0.00744965010097565,-0.0031706893761404,-0.00042200927141911,-0.0318195261239941,-0.0121341128517161,0.020223441340782,-0.00589103658931234
"524",-0.00301815664086058,-0.0128056805789916,0,-0.0101548220720116,0.0186055692104607,0.00811098345064942,0.00638163341002773,-0.00465935877560486,-0.0270507288807519,-0.0192592500730235
"525",0.0140468597463461,0.0335749242154362,0.0189800529655026,0.0298844060013372,-0.0238166495015676,-0.00861313643933992,-0.00380478975160181,0.0144684768567789,-0.00416473454141086,-0.0115811681446749
"526",-0.00489621814618457,-0.00996679689882896,0.00931310303833621,0.00736248385792337,-0.00349917820727563,-0.00508541302122334,-0.0235517804447692,-0.0151009712618817,0.00802530792330391,0.00560380148302553
"527",0.0148806887118385,0.0193884280870196,-0.00346026212824813,0.021066040603539,0.00087802964107242,0.00234246580077735,-0.0153190478581801,0.000426136260400556,0.0105405135680645,0.0222897741548633
"528",0.0284971936997176,0.0263350259342958,0.00578696637727605,0.050105145849882,-0.0031187094398385,-0.00605642010469987,0.0685198410060059,0.0400166604243888,-0.00588112497066828,0.00743300010297254
"529",0.00137948313437652,0.00819669748314023,-0.0184119031776862,-0.00521245043314911,0.00322616260060249,-0.00203019559650242,0.0136312762135702,0.012280439775505,-0.0141756452361044,-0.00541064938474589
"530",-0.0458091608483691,-0.0516082387529377,-0.0351701925139543,-0.0604594027971841,0.0217307510680642,0.0133888094524048,-0.0858804762646211,-0.0477155736678019,0.0213994451992754,-0.0128586343260043
"531",0.00589577536769315,0.00782711560853722,0.00486044247886053,0.0300299107326238,0.0129712408139402,0.007715361524542,0.0254097343965165,0.00127396463300911,0.0230573331455197,-0.00601204533501087
"532",0.000717673666239094,-0.00517782917522358,-0.00120912430729359,-0.00624725663229231,-0.00941587255756571,-0.000314072575491986,-0.014672380827933,-0.0029686143692097,0.00953512829629299,0.00151228372584122
"533",-0.0107575513702696,-0.0115239184020371,-0.0266345001386753,0.00502912911417641,-0.026613387070088,-0.00786915192880588,-0.0598943761641063,-0.0110587895803168,-0.00665444899977352,-0.018117878429032
"534",-0.0427743146115072,-0.0590450031312414,-0.0335821383168911,-0.0638033065048638,0.031148898297622,0.0168148047413228,-0.0630058789391671,-0.0692477051381304,0.03133434798484,-0.0558688131967552
"535",-0.00239843386080296,-0.00439636578487335,0.00772201503176984,-0.00712656203780304,-0.00852221318342394,-0.00728036036226987,0.00413233680190106,-0.0189467277820532,0.0152960402921751,-0.00597174427432889
"536",-0.0107553850224876,0,-0.0140484997550954,-0.0094215945379531,-0.0170011551236462,-0.00555299365071971,-0.0385333420007447,-0.0254350631064896,-0.0117635636461226,0.0245768480119914
"537",-0.00972134143437831,-0.012444478822203,-0.0129532888915989,-0.0253619967414218,0.0097160447306337,0.00284511370059737,0.0642021171086238,0,0.0211966802087298,-0.0111942597399849
"538",-0.0357787200410553,-0.0402441854369061,-0.0419948379312769,-0.0246284838657137,0.00923840552186683,0.000945481413687999,-0.0760512237017676,-0.0362497159070082,-0.0007157463993126,-0.00970331719433548
"539",0.0379099358951609,0.0427785787104047,0.0410959281557497,0.0547881079521131,-0.00104893276328366,-0.00377895047979848,0.082311082229541,0.0275828171062134,-0.0306968168209306,0.0190527660614423
"540",-0.00787292579733401,-0.0288383991466918,-0.026315825856707,-0.0171636005815947,-0.0115488714452602,-0.00906002610618528,-0.0252282398971784,-0.0278184197066988,-0.0166789923990607,0.0117521957846016
"541",-0.0162610049340659,-0.000836319340817071,-0.0121621530615085,-0.00873152239036867,-0.0105255037680188,-0.0025515148630465,-0.0423858360836766,0.0115462678349969,-0.000966226495625944,0.0211193055324381
"542",-0.0223490373416348,-0.00711601854770838,0.00820773646535011,-0.0157630223826939,-0.00575759566993328,-0.000852326800752978,-0.0152761021328355,0.0143918551043265,-0.0046206856785016,-0.0118925004637856
"543",-0.0450424733288872,-0.0619731691552545,-0.0352776777523777,-0.0607628199669272,0.016555304115581,0.010032281155832,-0.0700082282339526,-0.0631115802073938,-0.0183525537629025,-0.0502355994577631
"544",-0.007507090105352,-0.00898872498281489,-0.00281325088584661,0.0140425156845654,-0.00668107887827729,-0.00127025849709883,0.00384954279099126,0.00574421922035651,-0.0097877378203014,0.00661170746738571
"545",0.0236907651274381,0.0380955175253235,0.0267983816502342,0.0702272412047171,-0.00458093925356728,-0.00508980762934907,0.0264170421270775,0.0150569014703477,-0.0116615169739948,0.0350300751350248
"546",-0.0408474831282377,-0.0397555506647502,-0.0192306756524598,-0.0411275509791194,0.0278099166528811,0.0117234897011456,-0.0643423668903879,-0.0424550160522906,0.033711653752369,-0.00846112494133433
"547",0.00174407681853062,-0.00136507904616456,-0.00280130476958884,0.0168676771960092,-0.00666928925706245,-0.00474040892128957,-0.0146403144640638,-0.018696359685435,0.00326125672923716,0.0240000562089202
"548",-0.0117526750180763,-0.0241454751421872,-0.0351120623256836,-0.0194314513651546,-0.00585054570376242,0.000423882360256478,0.0211611802403537,-0.0446383543121378,-0.0186369160403412,-0.00572919525600046
"549",0.0596092227235359,0.0732958311515424,0.0509459928514622,0.0811986924254366,-0.0191991149049312,-0.00730063421279892,0.132275406070226,0.0717947017019889,-0.0268300872253504,-0.00261919038814651
"550",0.00651270638148271,0.00521976000176649,0.00415506550793765,0,0.0108206390048806,0.00714092292161728,-0.0171340858605374,0.0159494560754148,0.012253256322365,-0.0315125524628562
"551",0.0393718553714837,0.0359150411560176,-0.00137931839807426,0.0384442806527894,0.00476825363296185,0.00285643349788001,0.0788430016785733,0.0387228378153928,0.0210714747694298,0.0466376618266351
"552",0.00781481298292008,0.00167066022097373,0.00966844041865622,0.00559630996938365,-0.00503692358495644,-0.000738241853447619,-0.0212997739101057,0.0292195005415563,0.00219544461460908,-0.00880838321565069
"553",-0.00302303861451425,0.010425413380561,0.0177839218322078,0.000855976032455352,-0.0157685212656145,-0.00570216556801939,-0.0735460031601366,0.0234947393430689,-0.00547645107963468,0.0219551233768189
"554",0.0305831047434071,0.0222868204118025,0.034945997164531,0.0218134362162381,-0.00543964369864613,-0.00191190532542884,0.0745241457292958,0.032520199137718,-0.00837006580275113,0.0214833462568833
"555",0.0223844678784229,0.027048624499501,0.0233768045468781,0.0209290375167783,0.037887256183714,0.034262476994283,0.0516396592659167,0.0310332069066936,0.0338737779445382,0.0125188655265474
"556",-0.0123863668387461,0.00353781694901456,-0.00507617210753153,-0.00655960705274372,0.00124546835847927,-0.00339503489929327,-0.0569897354502732,-0.00628989639554345,0.0135353104967368,0.0207713816451687
"557",-0.0212939386649719,-0.011750800851671,-0.0216836107070738,-0.0136196298793877,-0.00555050558465697,0,-0.0744959854572932,-0.0134089416030865,-0.0080551353058852,0.0135659568000472
"558",0.0718293052844572,0.0729293315219599,0.0782268866185336,0.092468825143259,-0.00865990866973809,-0.00340650722606606,0.149897463839328,0.0411023221699049,-0.0161341389522017,0.021032562538039
"559",-0.0197035628568247,-0.0369417078753961,-0.0278114200244387,-0.0310228405025056,0.00951273718226897,-0.00145062877591873,-0.0714286960089736,0.00897265566973826,-0.0122719914797569,-0.0163857844833152
"560",0.0105462349620293,0.0149598875257109,0.0298508850389241,0.0150198483877579,-0.0134620057647171,-0.00601554065510512,0.0138824368975046,-0.00222385677988468,0.0113249701371623,-0.0152308792253397
"561",0.0203809503942434,0.0120936182666271,0.0108695191073438,0.0272585598330362,0.0115989035787281,0.00260873218213775,0.0248262467505305,0.0160430294353899,-0.000543629032062398,0.0173997215694346
"562",-0.0180488017035397,-0.0403286870552241,-0.016726608615658,-0.0295677541014017,0.00741844280599846,-0.000624595539683859,-0.0401212203910098,-0.00350896143993307,-0.0134885021211791,-0.0185273076455011
"563",-0.0345547799098918,-0.0412451482814767,-0.0388822266315727,-0.0515623802711396,0.00382552557272531,0.00427036086299704,-0.0548108747920982,-0.0528165710296815,-0.0078288563716209,-0.0363020355662409
"564",0.00926506427946427,0.0381492707765163,-0.00126400250735836,0.0218284540984717,0.00714584314253441,0.00176279544259939,0.0621609524420421,0.0250927538020804,0.00333402967323759,0.00452038323437498
"565",0.0193662849573104,0.0234559998223014,0.0291139055309106,0.0330511842062164,0.00912620416601184,0.00245080274539067,-0.00903375382939131,0.0117857262415813,0.00830748790770364,-0.00249996577856626
"566",0.0292379342235252,0.0469823957033566,0.0356704935993564,0.0542335140771402,-0.0122211834968753,-0.00652550345204006,0.0661913964691743,0.0640685085140178,-0.024497374761039,0.0385963742912467
"567",0.00994794323201154,0.00839127928834316,-0.00831372983027201,0.0122129360397343,-0.0204627287299588,-0.011467605853351,0.0895903111097722,0.00505255173874386,-0.0136262044946103,0.015444053609444
"568",-0.00783243302328673,-0.0188132787654252,-0.021557014885191,-0.0124312914598264,-0.00427537989528692,-0.00231992945322446,-0.0160350309364879,-0.0146624286546015,-0.0264870316925234,-0.0123573436304513
"569",-0.0233258890917654,-0.0265487574681377,-0.00611969440551852,-0.0229546366138192,0.00253737141683374,0.00253660219698815,-0.0752427880736043,-0.0153062721533518,0.0172393696694981,-0.0178056351805647
"570",0.010778355039732,0.0102271331876664,0.00738924269773378,0.0147784429468221,0.00885733752034068,0.00495543717699332,0.0209973348463426,0.0250428197890273,-0.00149869729072394,0.00734928855250017
"571",0.039742280963623,0.0217476343555281,0.0366746976402135,0.0436893343193479,-0.0125424128023297,-0.00587627072996744,0.119353803513115,0.0421230491946196,-0.00346383785401416,0.0145914913061271
"572",0.000233646412192146,0.0176143374297559,0.00235850442639096,0.0060821918771492,0.0091847469167945,0.00591100539797207,0.0127950412214739,0.00525496110358836,0.0181902333029831,0.00431451718146958
"573",-0.0172438137279178,-0.00937606032618865,-0.00941167861050918,-0.01600266528886,0.00522765282961957,0.00514103016017864,-0.0819565265236695,0.0072375579322892,-0.00580330015259334,-0.0181385200973956
"574",0.0106701261356326,0.0152895175206318,0.00475047864541556,0.0144560967036329,-0.00173362245922271,0.000939722519271324,0.0818633191509903,0.00518992843483002,0.00148789052920151,-0.00631979731497179
"575",0.0146627082816275,0.00609523333107087,0.00354583629139071,0.00855001267961852,-0.00791151157795555,-0.00396307278343089,0.0407693779588869,-0.00198576323009214,-0.0193143085714287,-0.00440312116309871
"576",0.00670557257347437,-0.00178197574612371,0.00471177244029852,-0.00706473416983433,-0.0109880628825159,-0.00806152736027466,0.0100284766365761,0.000795663666328439,-0.00687562071729675,-0.0073710074952722
"577",-0.0419154776349652,-0.0485540269664984,-0.0222745256484954,-0.0487370782439769,0.0151416949359304,0.00696657467068795,-0.107043062634595,-0.0588467973834165,0.0203003517918288,-0.0376237562217255
"578",0.0195375916108167,0.0228892970040477,0.011990299770273,0.0213162864983236,-0.00987949383290421,-0.00387841049567883,0.0913822802980839,0.0190115150145342,-0.000690028775964135,0.00360077366973188
"579",-0.00611398188799017,-0.0110050097956278,0.00355473753718316,-0.00842165624106905,-0.00606567845602368,-0.00242052515906344,-0.0337468815401942,-0.00373153378570878,0.00563929112256067,0.00153775748535745
"580",0.00981813582423774,0.0315279816118683,0.00590332878655841,0.0155094462833503,-0.000098121405818663,-0.000210628999157914,0.0415155106320142,0.022888214574041,0.0162509275435201,0.0133059086425964
"581",0.0151105718968949,0.0172600552926614,0.0152580217087714,0.0189092867261518,-0.0100405784867498,-0.00390387557184979,0.0528312859375843,-0.00325508033037558,0.0103603374878263,0.0151515687072972
"582",-0.0094623733433512,-0.0130787065921893,-0.00231208303730057,-0.0335475044158847,0.00427542425292637,0.00413067458453531,-0.056490408818912,-0.0191834296398533,-0.00791349745972469,-0.0248755890277783
"583",-0.0031454400232056,-0.00286526614973237,-0.0162227490289989,-0.00332375518410621,-0.0163366838186761,-0.00485289159795288,0.010828314863861,-0.00457782870016898,-0.0141557349925686,-0.00714296929139702
"584",0.0212694998201259,0.0312498184518768,0.00824550452871042,0.0526122363832138,-0.00885768564881717,-0.00540575188861447,0.0396973586545357,0.029264182055893,0.00660970940170924,0.0231244135623185
"585",0.00034270713781237,0.00452805573220783,-0.00584136490612641,0.0091516907554432,-0.00396034741993245,-0.0017050427031664,0,0.0125917017093071,-0.0120005091814669,0.00351577321474195
"586",0.00537666910095025,0.0124826563396991,0.0152762357080518,0.0146494468885043,-0.00688215884475063,-0.00321207600423057,-0.0339393827914609,-0.000401284618166686,-0.0036667813796305,0.0300301367672682
"587",0.0340198251722825,0.0410957564730448,0.0266203858535849,0.0690960306754882,0.00329462213324061,0.000965964919119378,0.0865744822691983,0.0389247823754435,0.0194364814066641,0.0194363296856011
"588",-0.00341085310824529,-0.0108551123597767,-0.0033821390310006,-0.00900330137930028,-0.00123148653974781,-0.000214379856005142,-0.0334870456555129,0.0023174958543013,-0.0043998082626332,-0.014299382269237
"589",0.0173341260105537,0.0216164014350007,0.0237554868049241,0.0171967488805047,-0.00236374507786419,0.000429388436324674,0.0334527468412311,0.0354525119361275,0.0146175750708215,0.0265957801542649
"590",-0.0138915291451164,-0.0179036660565645,-0.0232042583518292,-0.0248804959927689,-0.024412330978926,-0.00836827693681452,-0.0578037227563216,-0.00744340481339112,-0.00111680811797177,0.00188410047824861
"591",0.0233324279754263,0.0477293129321126,0.0407238420626104,0.0333662103585051,0.00242819618525081,0.00118976204453891,0.0677920012793778,0.0292470386261785,0.00603757812974992,0.024917674809716
"592",-0.0187135570133595,-0.0306863901602801,-0.00978260089241256,-0.0234252053371651,0.014219593111263,0.00940268815433365,-0.0293017210787871,-0.0280512397305789,-0.0032229494368875,-0.0082568156770203
"593",-0.00295970569852533,0.00979119342488621,0.00548830867399541,0.00713134550632044,0.00363451941352144,-0.000642996889104408,-0.0159815592378071,0,0.0112609541473752,0.0101757669694855
"594",-0.0251730607806818,-0.0303815854511892,-0.0185590311098247,-0.0366913393377341,0.0108653890665817,0.00460698584257657,-0.0679699105702724,-0.0431034368559238,0.00429987886328154,-0.0114468713857856
"595",0.00857074076773778,0.0103336281646251,0.00111262100187526,0.0143668312301752,0.00389034156858648,0.000106617987858826,0.0319457514263923,0.00940033560396691,-0.000658656302937932,0.00648449018123598
"596",-0.00816197173595179,-0.0131972745176756,0.00999989159014736,-0.00922262449113453,-0.000306278212637068,-0.00245254022783159,-0.0328325365425539,-0.00388045641813184,0.00571244650897995,-0.0253106155559778
"597",0.0284069855848639,0.0434637475695741,0.00880109754047487,0.055518569302579,-0.0155040054336747,-0.00587912290947401,0.0750075673725281,0.0268796567362333,-0.0129983829711071,0.0264399184207804
"598",-0.00120578447659569,0.012496131910384,-0.00654321094761701,0.0113383106443314,-0.00528378430035403,-0.00139839190652546,-0.0159396654566725,0.0170717748593929,0.00664008403452754,0
"599",-0.00669413784996564,0.00474686973860416,0.0131722505861878,0.00311459129915503,0.0105197355410278,0.00312282569493472,-0.0116137989952437,0.0104435564417544,0.0141820691972523,0.0160994686754468
"600",-0.0143631103036321,-0.00440958388486179,-0.0130009981802863,-0.0186278816249945,-0.0251497164572476,-0.0109476364814042,0.00185551047070032,-0.0103356158542205,0.0173441517615176,-0.00814846504239086
"601",-0.00213000709607347,0.00379638380271885,0.00329316974739213,0.00442908050624236,-0.0111012664207876,-0.00586119224983328,-0.0212964726717101,0.00522132722720281,0.00319663299300221,0.0146050497443448
"602",0.0256118593065882,0.0211158895302386,0.0328223884752272,0.0119684901516448,-0.0150752539179976,-0.00665989435302705,0.0517185800066202,0.0330241735984416,-0.00414232598741737,0.00224927486095283
"603",-0.0178526471865994,-0.0169754562151959,-0.0190675956234816,-0.0115157920022416,-0.0176953807758691,-0.0113198936148371,-0.0332831557252966,-0.0114940063430413,-0.00330636725029088,0.0044882691767838
"604",0.0139397409696762,0.0128727272727274,-0.00647942282279168,0.0308563820311019,0.0144779161564372,0.0052248420716372,0.0189207316880862,0.0148987119971011,0.00845372953837553,0.0183200938637791
"605",0.0177080151813718,0.0136392078933221,0.0184784346689937,0.0152720600741767,0.0258165389791545,0.0112786683091191,0.0273970270655473,0.0329390201545616,0.0207979524787341,0.0193066290542936
"606",0.0242084868524597,0.0284405294619645,0.0160084369464744,0.0421176824464831,-0.0295639077772476,-0.0163184775552861,0.0420740298056159,0.0183708017487589,-0.00488559266794986,0.027550648242207
"607",0.000843701613403747,0.00713624297744531,0.0010501739841422,-0.0144342441443809,0.0053792711837819,0.00334397037753353,-0.0147849291031554,0.0139551834302751,0.00658098798973183,0.00418930158616559
"608",-0.0126517291460362,-0.0345437643721963,-0.0220354005662382,-0.0354419805746249,0.00939038924601543,0.00611194877390542,-0.00230888608795765,-0.0184624493603156,-0.0202365813591056,-0.0333750258162775
"609",0.00939683596899554,0.00795101309547763,0.00751057965018953,0.0185238720032641,-0.0206614744199141,-0.0115969853034348,0.0295050987782302,0.00273523445752866,0.0192776074874437,0.0366854001460537
"610",0.000211587501936839,-0.0127428112442122,-0.0117146592778513,0.0020871461166434,-0.00762180399433199,-0.00994528127456851,-0.012644047452698,-0.0225097925762945,-0.0261873004410069,-0.00541225372086029
"611",-0.00412463088839776,-0.00522421933422745,0.00538802798117666,-0.0154715946819071,-0.00256007821805726,-0.00507855501556553,-0.00369963983917376,-0.000348864182597941,-0.00160069364636317,-0.00251151998290522
"612",0.00509754547644947,0.0120482801906954,0.00857450920258906,0.00181337094071843,-0.000111600124585998,0.00431003170549848,0.00114294681286253,0.0150087973672113,0.00288589146827478,0.00965169779847508
"613",-0.00253579295271356,0.00274714365105644,0.00106254597692756,0.0126696699129962,-0.0157368200272754,-0.00598631789535753,-0.0191157889924932,0.00447081925594373,0.000319716501764544,-0.00374059749461575
"614",0.0044494691676209,0.0167430061940017,0.0169850809636907,0.0214476559800185,0.0111122114770861,0.00681817092256654,-0.0186155737201706,0.00581946390396992,-0.00170470912311205,0.00917814283389506
"615",0.0027419183141344,-0.00508995447514538,-0.00104369099526413,-0.0160397160343811,0.00897205224099262,0.00530490441445375,0.028156617931,0.00646686635596616,-0.0163286984950489,-0.0140553730163712
"616",-0.0229282423995107,-0.0373158054853783,-0.0177639506710081,-0.0358624518516732,0.00900248931906877,0.00449056932646075,-0.044969580165785,-0.0246868745023227,-0.0116089836521425,-0.0192872499722414
"617",-0.0135628928382009,-0.0128163057866972,-0.0106385217741978,-0.0150630173827433,0.017404932951526,0.00558896443901835,-0.0141865959633307,-0.0149099153110465,0.00911088933284065,-0.00384783372232922
"618",-0.000982115809816109,0.00316643518140158,0.0118283538703108,-0.0112359219195047,-0.00562959776415406,-0.0026679399412487,-0.0140844200075098,0.00457599349010462,0.00456867181551179,0.00300442766130105
"619",0.00731813370392476,-0.00315644051710029,-0.00850161205181399,-0.00284086084836488,-0.015135194911517,-0.0121478715038156,0.00496893375764529,-0.00455514915721467,-0.00801296173281996,0.00128359132876055
"620",0.00368594146468926,0.014566002649028,0.0160769754933441,0.00506485644495047,0.0137087396644284,0.00462545769220379,0.0108156746299546,0.00997142033827703,0.00316560415712686,-0.0085468920092806
"621",-0.0299870077516331,-0.0362213516657621,-0.0221519384193041,-0.0362205800492651,0.00970703644421356,0.00539024921983411,-0.0510548075464354,-0.0278561352190982,-0.0147987047921936,-0.033620804004005
"622",0.000784030939245062,0.0201985583005344,0.00650773437722907,0.00649008542088936,0.0117728044662815,0.0032398282385977,0.00869855551347198,0.00652895382691088,0.00419700680144675,0.017395175235059
"623",0.00861801809143414,0.00194748543883749,0.00215504759335583,0.0219314305260894,-0.0100342548242475,-0.00378599430191495,0.0164382477776746,0.00504490016803527,0.00582928961349061,-0.000438398234711701
"624",0.0217483801909122,0.012957644286973,0.0236560879763297,0.0297886119006658,0.0183328206412994,0.0125170069543405,0.0159489913440176,0.0340627048943116,0.00940405717017123,0.0087719456635289
"625",-0.00260576187080441,-0.00319788490315143,0.00315134445110088,0.00528782298336794,0.00169391877568748,0.00132447583767115,0.00879117444155297,0.00970826623312826,-0.000216628755641324,-0.00826089106396555
"626",0.00936362803377566,0.0112287032021163,-0.00523565775143053,0.00742585637353543,0.00148002769211941,0.00209391830243555,0.00248949057573955,0.0058380889688241,-0.00270885250071673,0.00964489652745826
"627",-0.00809048770088339,-0.00444190452318438,-0.0073682923517534,-0.0101352269403754,-0.00168910810112877,-0.00263993412912311,0.00651964456909337,-0.019119171660954,-0.00934377434437439,-0.0178027572355389
"628",0.0041328044075406,0.0152966223980513,0.0116649020782458,0.0183055649229116,-0.00198399088608381,-0.000640267194878752,0.00987081123302924,0.015662969882217,0.0132704430796227,-0.00397881616864659
"629",-0.0272932831904782,-0.031073519988789,-0.0220123790113054,-0.0274220760508256,0.00233914903661336,0.00331933253576677,-0.0455102655248347,-0.0215895785511684,-0.0123389870368978,-0.0221926019969989
"630",-0.000111425020806188,-0.00161946047361972,0.0064307811094797,-0.00219271449213732,-0.00190904378237911,0.000661619580328399,0.0208001546295749,0.00910628971919047,-0.00536984109589045,-0.0299592023076115
"631",-0.0193769300950973,-0.0295264889243423,-0.0106498020051367,-0.023548164038156,0.00669380546900022,0.00396896179214701,-0.0369907500883468,-0.035751203876707,-0.000550936523778467,-0.0159100812892855
"632",-0.000680926954879979,-0.00668672215780741,0,-0.0115755205016084,0.0184696425289184,0.0115277866271191,-0.00976547727515364,-0.0104391386127212,-0.0158747879602555,-0.0123634141565601
"633",0.00193189233676261,0.0151464393770202,0,0.0178919596395444,-0.0119174395486707,-0.00586121351995872,-0.0161078138779669,0.0080029566911759,0.00268852927148622,0.00625904125719567
"634",-0.00238181701633744,-0.00795782750925911,-0.0107642804658418,-0.0118248687052079,0.00922943311873037,0.00622337374769222,-0.00167082645036265,0.00360872979664673,0.000782035509282908,-0.00765554569948457
"635",0.0243289863620715,0.0257355925945031,0.00217637967831141,0.0071152019509757,-0.00561202520000548,-0.00358103620737416,0.0394916770141158,0.00898968173589965,0.00680955555236551,0.00530393685595221
"636",0.00566083206758461,0.00260675514536435,0,0.0109184971414915,-0.0166160572343321,-0.00664264491209954,0.0115902232957015,0.0242335246641401,0.00687433181340857,0
"637",0.0292459899097368,0.0425737789418663,0.0108577155324761,0.053684750469625,-0.0257172359058234,-0.0129352635864348,0.0343733017388019,0.0208767133348,0.0157471647560217,0.0263786816745606
"638",-0.00160833809706484,0.0109102281411158,-0.00429665481650587,0.00180886310141548,0.0107982294024078,0.00599757305513515,0.0129229803112305,0.0248805901368225,-0.00281867959277282,0.00233656119252856
"639",0.0109548146306602,-0.0037003175408894,0,0.0102318167549371,-0.0154308696866046,-0.00673495512546896,-0.0233902249448401,-0.00897866281286563,-0.000543629032062398,0.014918402839005
"640",0.0106236041573671,0.0194984783436423,0.0129453294838178,0.0357465642564436,0.00526072645142572,0.00366841666801743,0.0323484941822123,0.0218116551800343,0.0146850756010006,0.0165364813130622
"641",0.00462528900820613,0.0045540346117654,0.00851968260912539,-0.00287642414067057,0.0199522059309845,0.0111846611168576,-0.00210915265068901,-0.00426880186260048,-0.00160808320763384,-0.00361499950632049
"642",-0.000209104606818888,0.00392841650068765,0.0116155038098773,-0.00230751792844763,-0.00897930318343088,-0.00591426707907461,0.000906094947973113,-0.0042879515976233,0.00332873413493195,0.00544224272584604
"643",0.0220826357301411,0.0174596633300323,0.00417534094337246,0.0283316774661435,-0.018336146738378,-0.00969462685249867,0.0346904151948437,0.021530442234643,-0.00192636982178152,0.0207486147016711
"644",0.00409560312441481,0.00739618934488884,0.00519731199590012,-0.00477909177475877,0.00483448938292264,0.0021136474981942,0.00874653331469077,0.000648506884140865,0.00160842801611771,0.000883861571832734
"645",0.00295756607710063,0.00146845826222886,-0.00206841051794748,0.0087570661757812,-0.0114816324576174,-0.00466206265794999,0.018786176417863,-0.0116657374526016,0.00321159391021975,0.00397354664689109
"646",-0.00467763484778416,-0.0058649378637502,-0.00103600848906893,-0.00448042004366622,0.00884944641980367,0.00200679634193635,-0.00397165930965304,0.00557387862200387,-0.0170739303924227,-0.0109938289580486
"647",-0.00245148708685394,-0.00973465812086149,0.00726174861434736,-0.0225034852233456,0.00548258753749109,0.000668098516498183,-0.0142411137411822,-0.0091296608952266,-0.00987953523092455,-0.0257892071251772
"648",0.0104456003859141,0.0196605426054086,0.0113280049988884,0.0247480245631391,0.0141765484394099,0.00400462428847348,0.0349609879016124,0.0164528061807874,0.00460532909885947,0.0310360066831867
"649",0.00141864548180437,0.0169442488420435,0.0050919179041542,0.0047737576617326,0.0194619549912336,0.0100817346171709,0.000837457420632903,0.0213665087663568,0.018882284908897,0.0199203653748934
"650",0.0164965549875562,0.0264291268764996,0.0172237425975421,0.0374509964178138,-0.0151542197140634,-0.0106265531616068,0.0198048781313818,0.0288430339051875,0.00557048753230815,0.0282116866853799
"651",0.00258812567293321,-0.00335863531447622,-0.000995854171498833,-0.00915930392158615,-0.00795231515697181,-0.00289040265222906,0.0475930795167487,0.00462117411591945,0.0086289227028149,0.00042220018779604
"652",-0.00287937143546002,0.000842430501221791,-0.00697894037780922,-0.00842839661624617,-0.0149478594004192,-0.00568746883547167,0.0404698969679287,0.00275993898275106,0.0010561787072243,0.010548596042903
"653",-0.0051787576720016,-0.00841756143466388,-0.00100409254727574,-0.008225834683106,0.00340832639220867,0,-0.0062734810911641,0.00152882313173341,-0.00189914540936009,-0.0229646233327346
"654",0.0131139906986262,0.00028322804621661,-0.00402016697539243,0.00995282393036701,-0.00832874514623638,-0.00661609595169543,0.0464646940022695,0.000915916095461045,-0.0089851798939784,-0.004700702637916
"655",-0.0020748626234246,-0.00735491814626366,0,-0.011223644619402,0.0124879571932786,0.00643439693256975,-0.0197879475607671,-0.00274551432317161,-0.00874666666666657,-0.000429451290466343
"656",-0.0124761998790921,-0.0108293844342887,0,-0.0188262478295225,0.0115695654080572,0.00695491547572291,-0.0295418414739443,-0.017130468997643,-0.00150649951576454,-0.0150343792638081
"657",0.0107291486941588,0.0146930908579643,0.00504555270220308,0.00902970954244475,-0.0106817357642202,-0.0027847028556871,0.00659562339166753,0.0289448400765642,0.00172428061510632,0.00523324715238638
"658",0.00763842377997337,0.0167519213098231,0.00903617338360596,0.0173375679597039,0.0141774990404928,0.00781941002075892,0.00478845276003059,0.00574694585403557,0.00828406696990003,0.013449063960312
"659",-0.00767951278374268,-0.00949468146194876,0.00397971923502549,-0.0181417304181964,0.00387202746875759,0.00310383746780762,-0.00902976219455265,0.00330842924536001,-0.00768246897479219,-0.0282533912361369
"660",-0.0246053530015597,-0.0352410930620359,-0.0277500335805814,-0.0391937306096767,0.0147833655931289,0.00685030599328496,-0.0501135216875052,-0.0344723403676045,-0.0149462258064517,-0.0149779951796416
"661",0.00793406524383444,0.0187025014981625,0.00815486614984073,0.0218531594896698,-0.00580618759333151,-0.00351125649881279,0.0122569533029182,0.0229741181348635,0.00491209469586185,0.0196779575566206
"662",0.00877971148232093,0.00975343104414761,0.00303326663355064,0.00256620620653858,0.0082819588309635,0.00374430628317879,-0.00737061161619068,-0.0145676040132027,0.0051053770390046,0.00701749333334312
"663",0.0103041341299519,0.00909078511411243,0.0120967964044865,0.0173492989075921,0.00821338339783861,0.00263313188979653,0.0405727714237927,0.0163224960056281,-0.00280992113703582,-0.00827519375240693
"664",0.0196059597313285,0.0295607828145847,0.0109562397855059,0.0150966908485208,-0.0205762422291864,-0.0101774748481626,0.0221711958087694,0.0148488450663045,0.0149561617521241,0.00746599767470402
"665",-0.0000969899862699464,-0.00136719308301847,-0.00197027029078334,0.00440624519225308,0.0181294586262037,0.00619135680720806,-0.00573408614867843,0.0050760752498975,-0.0139883179073504,0.00174365530253318
"666",0.001942200151686,0.00766706451779364,0.00789717024698278,-0.00219345768375312,0.00565611792724385,0.00263711732048244,0.0110331617435824,0.00950702971359174,0.00454847323146956,-0.0143603410888363
"667",0.0000973694277006665,-0.00407590667422475,0.000979506746570991,-0.00302300780725606,0.00458345474817246,0.0013150418546457,0.00446420976226469,0.00176574016079001,0.000323404477718725,-0.00264897051125457
"668",0.00222931960256423,0.00818536300835015,0.00293541102386485,-0.00192937431139595,-0.00394055447918573,-0.00273627305083168,0.00790129643016391,0.00793193320529606,0.00431082008502193,0.00841077740029217
"669",-0.000193730003362425,-0.000812102863980368,-0.000975771610715048,-0.00524710502051395,0.00458037880239415,0.00230484058933444,0.00661464546468449,-0.000583240453737921,0.00729693084457694,-0.00219496822668053
"670",-0.0088989856125119,-0.00622961759311302,-0.00195295363132586,-0.0197113994981231,0.000932189509642134,0.0029558939458012,-0.0124122360433074,-0.00670747979142272,-0.0050069349630254,-0.0272766279455596
"671",-0.0220577519651171,-0.0283453951371349,-0.0146772304183271,-0.018974692046149,-0.00241995834804676,0.00259493100505193,-0.0510102982792519,-0.0284788199646797,0.0053533189431838,-0.0153776794646028
"672",-0.00379234183437638,-0.00364670572068304,0.00297937371031765,0.0106815133378937,0.0145750091777859,0.00545995953316525,-0.019735186925022,0.00604388405672762,0.0243876459129362,0.00229675452761691
"673",0.00831500251248851,0.00760143377014755,-0.00297052341096116,0.0199940523510902,-0.00615617033065674,-0.00358422613411991,0.0177483794188831,0.0156203245314357,0.0132030041957998,-0.00504131910971206
"674",0.0140092541952797,0.019279220413122,-0.00198580436463025,0.0193224019987293,-0.0170346799539386,-0.00599416217843662,0.0119731815711726,0.020112127142611,0.000718243389270068,-0.0041454986395717
"675",0.00862178915754797,0.0249450519991163,0.00895510361875784,0.0206043379743701,-0.00703812580756336,-0.00230218082409051,0.0321500498561889,0.0171067443297406,-0.00102531529811656,0.0185013728514223
"676",0.00767470589629138,0.0117679180405248,0.00394475011743478,0.00538362363573519,-0.0011628487889398,0.000878464516968602,0.0201842674436332,0.0188141451763855,-0.00359230216565753,0.00408723115819432
"677",0.0102189454472024,0.0113665318759413,0.0117877212903552,0.0131190781660004,0.0184255990187716,0.00746669307203129,0.0141671244184562,0.012590749108212,0.00638643373740355,0.00542728758512201
"678",-0.000190897536344603,-0.00313618129195747,-0.000970947949067047,0.000528386987340035,0.00551167112748385,0.00294359977775205,-0.00313123452955755,-0.004420897483848,0.0110542685072959,-0.0130453034291789
"679",0.00486790877760934,0.0049816151159745,-0.00388713115461448,-0.00369734975239921,-0.00992802121098513,-0.00586886015649657,0.0287514326674356,0.00471832954478302,-0.00830127564589267,-0.00546948107058731
"680",0.0041793667254566,0.00391313821433692,-0.0078050367771455,0.0119297555320337,-0.00511729988838772,-0.00207650424965877,0.0176134531103984,0.00414333115109122,0.00959578409142292,0.0233729683713699
"681",0.0151341789721255,0.01845131990029,0.00491659134810529,0.0251507325392029,0.00178483990161515,-0.000766784935001819,0.0390033517035953,0.0198076366020228,0.0102123557085469,0.0129871590421937
"682",-0.00149079322446444,-0.000765614872204057,-0.00978460602454767,-0.00536693180513825,0.0125757649301854,0.00493264784908964,-0.004886693772303,-0.012139265808443,-0.00570521446480976,0.000441898573175337
"683",0.000637270904344955,0.000766201487458096,0.00494040923826611,0.00282636873396935,-0.00890093814746518,-0.00534488766862506,-0.000223377979118311,0.00607254916678235,-0.00674449392971577,-0.00883775159514855
"684",-0.00252980127163394,-0.00918590437528521,-0.00983280101431072,-0.00871129903167556,0.00229714971855888,-0.000658132529345878,-0.0158517241185356,-0.0148152447254841,-0.00314175540978534,-0.0218456740229847
"685",0.00582419307617354,0.0113310803960809,0.0129097298602132,0.0152495394003553,0.00208398426730549,0.00263365171023144,0.030923033764654,0.0158731710514459,0.0133183914872064,0.0164083024803074
"686",-0.00831209284870205,-0.00789414130933264,-0.0107844930417961,-0.0150204839387195,0.00301531553949541,0.00218953683441381,-0.0335254314258702,-0.0175438141604158,-0.00842777181554688,-0.022421542462665
"687",-0.0110190265411151,-0.0202769244749859,0.000991392865694163,-0.019643433421625,0.00290250300202688,0.00273053313165161,-0.0330809088663014,-0.0181360343415252,-0.0129515225548613,-0.0128440036923365
"688",-0.00533295113935173,-0.00445371112263848,-0.00792086361732469,0.00421848326622731,0.0127132332826456,0.00402948806501957,-0.000712707914835242,-0.000852737897565126,-0.00563816487017432,-0.00789966405563647
"689",0.0179037845404419,0.0142100987397389,0.0079841046211353,0.0128643038084824,0.00877706838139258,0.00173550046123694,0.0389920029874757,0.0145053468742784,0.000515494845360953,0.00889941747812428
"690",-0.0030100056609822,-0.00155659151462584,-0.020792244822759,0.00233244173301084,-0.000910263462922334,-0.000432227702484633,-0.0167050433486239,-0.00616788418690983,0.00391547643744028,-0.00371406505878014
"691",-0.00386798983246406,0.00155901826923488,0.00505566579263661,0.00620674983074565,-0.000912046604159,0.000757446568553366,-0.00698140161024019,-0.00310279932841606,0.0145745458277737,0.0279589470361863
"692",-0.0248131099037427,-0.0298388404040978,-0.0251507825244963,-0.0272424636045513,0.0136960380843807,0.00752317189365703,-0.0424185968466496,-0.0200906580851326,-0.00971167445041321,-0.00634633504819593
"693",-0.00466134428806775,-0.00909338954099448,-0.0134159905860438,0.000264074174533002,-0.00692091419152852,-0.000430631615737531,-0.00978969044323663,0.00664169772813961,0.00490350398307782,-0.0100365005487431
"694",0.0149279412617036,0.0145747969106216,0.00836812098873496,0.0232438793497647,0.000100977830164162,-0.000107295488177006,0.0269403031656836,0.00114785155615071,0.014740235394727,0.0322580997056205
"695",0.014324320136516,0.0188883307492542,0.0114107307386211,0.0165204393738339,-0.00989665597722611,-0.00323492315502194,0.000240777516976598,0.015758791195704,0.0246443498296935,-0.0120535907304756
"696",0.00274866581695199,-0.00261130502726847,0.00923101545488092,-0.00101608207409465,0.0117296296424301,0.00638142471274983,-0.00312801510203053,0.0146686929189728,0.000782186163298615,0.00180756951475836
"697",0.00765603206245302,0.0172777482540289,0.0111788032269,0.0122015109906166,-0.010484461123453,-0.00365426840318972,0.0188270543083608,0.00917448729638726,0.0125048650595461,0.0198466927695415
"698",0.00609695329106796,-0.00643326595336091,0,0.000753091879029499,-0.0229242741811129,-0.00959944197491092,0.00971327777546938,-0.00247938580543972,-0.00771905642337956,0.00398048486315061
"699",0.00391584857621052,0.00880580541985432,0.00200999345977126,0.00828144591455926,0.00156456745400013,0.00294064974078179,-0.00164210485599003,0.00386614076596326,0.00700118658114302,0.0202642210679891
"700",-0.00204339328421332,0.00231078562261655,-0.00501521819140127,0.00174210257046825,0.0052051039980896,0.00228081067346864,-0.0150415524862664,-0.00687742745501507,0.00675940530628449,0.0112263661355538
"701",0.0172155127981954,0.0217723039058695,0.0110888955878266,0.0322978670423155,-0.0148110791017653,-0.00682665580341768,0.0367454713521063,0.0340719651153352,-0.000767331656103321,0.00768576514257147
"702",0.00365967183887728,0.00777137567086816,-0.00498521683659958,-0.00553534358248786,-0.00462599771891103,-0.00327223273562105,-0.00759509052085838,-0.00482190239171854,-0.0126703685928202,0.0101693954337263
"703",-0.00747429750518114,-0.0121890052839517,-0.0180359853848754,-0.0137947541861995,0.0081324335077011,0.00459629560550279,-0.0271337189854719,-0.01561220756091,0.00311101494156141,0.00251683053248986
"704",0.00826541611181963,0.0151097083565117,0.0163267417785635,0.0191411915039492,0.00785732821471874,0.00152597018723988,0.0231230447663986,0.0210555442424927,0.0101764198488079,0.0142258758004092
"705",-0.00528287734108013,-0.00297726776403795,-0.00301227764182721,-0.0132437098697402,0.00540613676919599,0.00228403761481943,-0.0186391875910848,0.00107083535436314,-0.00777132281191617,-0.00618816184932824
"706",-0.00897351084053766,-0.00273690398970239,-0.00302092782753727,-0.00536833995013641,-0.00599685723941012,-0.00227883267527129,-0.00783477271466815,-0.00642032914935131,0.00319089157205354,0.0211707498222049
"707",0.0101632051268417,0.00998034364525813,0.00201990351900139,0.00834156076628534,-0.00488889531812364,-0.00293702053571188,0.022493165859518,0.0123852822791561,0.00163853493975918,0.00812996973268176
"708",-0.0114332544687277,-0.0170456360238717,-0.0231852103912061,-0.00827255474816102,-0.00752553549508495,-0.00490952234945652,-0.0109990006156827,-0.0249995815358321,-0.00413779838602391,-0.00362906586020384
"709",-0.0108252377365761,-0.016084502316638,-0.00309611871524207,-0.0125121265274075,-0.0129542628319269,-0.00570152560510651,-0.0061523323906757,-0.0155487746788936,-0.0157502853560786,-0.0182111281800219
"710",-0.00458314784904623,-0.00740721872870598,-0.00414073196865161,-0.0173914433923393,0.0136571283704612,0.00860047185200208,-0.0152381335759313,-0.0135768947183448,-0.0000982034154898281,-0.00700753571954482
"711",-0.0188872453365144,-0.0270201488286953,-0.0103951206115573,-0.0457647877665985,0.00473696953070446,0.00306177423862675,-0.0418281769334973,-0.0410112900929821,-0.010996514698017,-0.0257368123829955
"712",0.0214533458796982,0.0330600053825492,0.0157562204190962,0.0442501152441608,-0.0108952759512797,-0.00479580517090417,0.0431491131273385,0.0330991434503654,0.0194579464074871,0.0311036398292528
"713",-0.028973090645508,-0.0358420592715268,-0.0124093514906507,-0.0466884769806521,0.0145109565185155,0.00744696342103524,-0.0191096457577771,-0.0221149154972435,-0.00155811663145167,-0.0252065640847321
"714",0.00733877257497872,0.00743464539861649,0.00942402136810183,0.0149054477477075,-0.00441980906114559,-0.00263137827656457,0.00147966110496989,0.0127573862562995,0.0138495856222527,0.0173801378940006
"715",0.00316354425562637,-0.0076435979755175,-0.00103729973616662,0.00157333410420279,-0.00999498343554772,-0.00230791575021083,0.0142819738093314,-0.00314924948138284,0.0241462440831046,0.0141666878942486
"716",0.00257992349663549,0.0143424192499124,-0.00207666066887169,0.0185915732992101,-0.00913951740568941,-0.00275389747753851,-0.0179653388378295,0.0103385067571848,0.00601163823043049,-0.000821681464220014
"717",0.0183950946730784,0.0172823095125509,0.00728395024136286,0.0205652005487429,0,0.000220826020877585,0.0207664307650408,0.00682203455995634,-0.00112040151485349,-0.00534540630864588
"718",0.00262037662967018,0.00205912973728162,-0.00619835724084505,-0.00125928305732936,0.00096505024641913,0.00298186379681864,-0.0154999443901298,-0.000564389758837103,0.00420636555786991,-0.0177759529768661
"719",0.0227762556047673,0.0300538435681008,0.0114344526480512,0.0368221944536182,0.00117902914614865,0.00044086298048418,0.0469862981206777,0.0364406018918813,0.00707439262775766,0.0164141340305319
"720",0.000182397527914935,-0.00274301196358506,-0.00719424151345538,-0.00462196310710272,-0.00181978030158347,0.000769945657436599,-0.0049344258952021,-0.015262794232761,0.00184857192257004,-0.00496887633467813
"721",0.00510997286915305,0.00175047938432438,-0.00103549209428044,0.00855348285265989,0.00418165518369507,0.00286032984507711,0.0184180635243791,0.0102403530961106,0.0111633823338257,0.00665829530987594
"722",-0.010167998905565,-0.0107340714871594,-0.0165800654911334,-0.022292195802544,-0.00181483992578324,0.000328827587905867,-0.0118246105155654,-0.0167122701253035,-0.0126824728591692,-0.0148822347476368
"723",0.00541130163961046,0.0126166453393388,0.00948379370248875,0.0171005370607804,0.00459919825606714,0.000767222892268604,0.0133736890389573,0.0189471304808817,0.0141391647180407,-0.000839266802493133
"724",0.0145046110026024,0.0174437288675633,0.00939435348884454,0.0250971854385653,0.0117124821272145,0.00536803602370162,0.0226904945551192,0.00929708276509644,0.0172225171719067,0.0289794580824827
"725",0.00116896859135851,-0.00612303583242113,-0.0113752079881788,-0.00356552999981974,0.00536669138792245,0.00217946626257137,-0.0142628151645405,-0.00623157479732894,0.00304581213954513,0.00489801833895021
"726",-0.000628863722804796,0.00073932218879369,-0.0104599872598395,-0.00787203196786046,-0.00586170155018462,-0.00250072968389514,0.0165363463926529,-0.00736080422703589,0.00250066086897682,0.000812252937989699
"727",-0.0130312552189449,-0.0177299464841264,-0.02325622501556,-0.0185142366203377,0.00179034883843987,0.00119949856740376,-0.0198823734761758,-0.0192254726709368,0.000445461024498828,-0.0142044773407461
"728",-0.00355138381736164,-0.0127847470865099,0.00757594901898395,-0.00416452793801603,-0.000210592505028195,-0.000108814183615746,-0.00760738073422873,-0.00588076727789288,0.00569901142389106,-0.00123505925958234
"729",0.0127024069166333,0.0210762929531372,0.010741123885309,0.0209103644065884,-0.00126149677491449,-0.00141603501596443,0.0113823334054268,0.00957751201531498,0.0119532404470826,0.00453423541191289
"730",0.00153392013153453,0,-0.0127524119128748,-0.00554222210270483,0.00631632176403296,0.00512470062013826,-0.0146992010466387,-0.00809140213345405,0.00384987309607254,-0.0114896742436308
"731",0.00351403670957784,0.0126835501995437,0.0172225594736901,0.0116306608233663,0.00460191596572845,0.00336334157721896,0.00396255158392678,0.00759482543675039,0.0164734589957258,0.0240763949254048
"732",-0.0162505879255606,-0.0348723245560241,-0.00846559305156758,-0.0388022076732638,0.00374856222162467,0.00454057858676449,-0.0283258862355967,-0.0304300190963304,-0.0133768218133213,-0.0113497883869876
"733",0.00337640616756696,0.000763472004964738,0.0202777269058381,0.00971808427980503,0.00238610055690591,0.00161414535114712,0.0375150561833937,0.0129570326426467,0.00504085703182455,0.0110701708064096
"734",0.0123705854334124,0.0218658752442302,0.0345187450426516,0.0286281547440184,-0.0111396099899114,-0.00551355359412553,0.0128970484771178,0.0264356230563372,0.0150466794798225,0.00729925362220607
"735",-0.000449448920629814,0.00273731467930949,-0.00404422468212806,0.00407838843614772,0.000839675163207598,-0.00205761891005274,0.0147797223291777,0.00138471810012808,0.0153348359686873,-0.00684387248095841
"736",-0.0078202284468103,-0.00719598183277059,0.0142129157265043,-0.00931904051266641,-0.0103852037288533,-0.00466654801146738,-0.00851481378411645,-0.0094027003021202,-0.00402754656821624,-0.000810606791958768
"737",0.00570748686077227,-0.00025003185989636,0,0.00916544031363786,-0.0105991584108416,-0.00741342288278346,0.0268928519723111,-0.00111658054571173,-0.0417017449461267,-0.00811360440726594
"738",-0.00153129523055395,-0.00599985832683991,-0.00800793234266906,-0.00860411680867479,0.0012850029936613,0.00274577442544,-0.0173856671244861,-0.00475153451067301,-0.00562636483516488,-0.00899800029003262
"739",-0.01109676178721,-0.0223844861671086,0.00302723520392134,-0.0185629451878319,0.00149736916577781,0.00350528527484784,-0.00604690800554686,-0.0235885177020387,-0.0190964899735082,-0.00990506872576724
"740",0.00374059768153168,-0.00128640017438386,0.00301812874876073,0.00614090834104219,-0.00459340174250733,-0.00196443630700649,-0.00135203402471529,0.0115039347319714,-0.000991446624374337,-0.0125052544077175
"741",0.00563512496241869,0.00154578902614144,-0.0080241454522888,0.00585946516114455,-0.0114848248402474,-0.00339075104881292,-0.00293339004330084,-0.00625536496835288,-0.000180404192724803,-0.00548755975720583
"742",0.00424774361101354,0.00360055491337996,0.00606686537217938,0.00364082102032159,-0.000107420686185189,-0.00493911196736574,0.0144834693773559,-0.00457776152109279,-0.0135354629128316,0.00509348414873867
"743",0.00684044686169316,0.011276121815265,0.0010051017624646,0.00677151100111772,0.00119411720096863,0,0.019406340372861,0.00919794129661811,0.00841564215148205,0.00548978970308478
"744",-0.0046483766105182,-0.0114036964814057,-0.00803229069056355,-0.0103291803713332,-0.00444731983500557,-0.00319815859165262,-0.00919060960755402,-0.00882942382109908,-0.000272124460669931,-0.00461984469599885
"745",0.00152696590694146,0.0110226755416358,0.0151822270405377,0.00582533183222145,-0.00119813881257957,0,0.00596307448220701,0.00373593015168594,0.0125215226614783,0.01729955854448
"746",-0.0120159510814914,-0.0268760976889071,-0.0139582082251046,-0.0287162898261986,0.016470666001797,0.00885187644292174,-0.00636646565242061,-0.0160323487157311,-0.0380858513517646,-0.0153464185073455
"747",0.00565729642148849,0.000260722429418436,-0.00202215762811997,0.00273278896551399,-0.00429215367489344,-0.0049354501230785,0.00773323588175723,-0.00212822157934023,0.0149990782559746,0.00421237281712639
"748",0.0101622525960308,0.00763780300276107,-0.00303941280534026,-0.00123869010967081,-0.0177828134641288,-0.0102498824654045,0.0120583416163287,0.00207335958079025,-0.0183570450213046,-0.00964764890606939
"749",0.00359346923239556,0.00833553551013644,0.00799830651871658,0.0100779708155554,-0.00559505651446646,-0.00445489127135912,0.0106155221694304,-0.00443373581209583,-0.00729311848414538,0.00720032777982405
"750",0.00196851413048615,0.0105915365175555,0.00305167212341728,0.00990332521589377,0.000220369739873494,-0.000447346905472434,0.0112892213455629,0.0142519271962041,0.00357921265101657,0.0176619629297825
"751",0.00473483295384769,0.00255634721602371,0.00709964506426597,0.0100518716671478,-0.0103699967021181,-0.00358120272446805,0.0126423605084147,0.0014634419925037,0.0169873106432479,0.00578508727199134
"752",0.00213337111737921,0.00484429566739308,-0.00402826787729549,0.0033979196641114,-0.0027862418455088,-0.00269535520259812,0.00359673484372514,0.00555394758672945,0.00175343298492603,0.017666362905564
"753",-0.00141983152298331,-0.00126843914477814,0.00404456045023505,-0.00358100434854436,0.00659539987442836,0.00264041201706777,-0.0143370729664545,0.00784875557876985,-0.00994935025473931,-0.00201862644316708
"754",-0.000355041573280257,-0.00152457342896717,-0.0110776547102747,0.00437124509534681,0.00657554919793157,0.00179993696680536,0.00171197897015296,0.00490323417619609,-0.00502466730227336,-0.00121349249101033
"755",-0.00959812640767288,-0.00865127133810706,-0.00814693367697283,0.00338481066215368,-0.00476059340816171,-0.00482983128298509,-0.0194322572986348,0.00143529063504744,0.00355370803329258,-0.0028351171688914
"756",0.0169596229343509,0.0266936689765154,0.0256675298040019,0.0291567295534378,-0.000890013434736159,0.00248356966241348,-0.00239535930243706,0.0214962448953113,0.0232038490952167,0.0251827673620635
"757",0.00264730435001992,0.00100030259563044,0.00600597923069568,0.007258158355123,0.00645833041423516,0.00439063115185756,0.00240111082558925,0.0103816731612201,-0.000910801432309705,0.00118857325538912
"758",0.000703985048407851,0.00124875372646227,0.00398017019980768,0.00209186783605908,-0.013387128763373,-0.00403576756098156,-0.000435552277922913,-0.00527642601035316,0.0164995902415568,0.0178076370356166
"759",0.00422149447456843,-0.003242594574143,-0.00891972633432381,-0.005799051667987,0.00168249241295126,0,0.00893224228698308,-0.00669983668920016,-0.00618780367343197,-0.0124417099344923
"760",0.00332732327188356,0.0080078658619529,0.0120000643926972,0.00793264076632028,-0.000447962316687867,0.00123893025658561,-0.00669409528177012,0.00533953857256031,0.00496303013896404,-0.000787390854466552
"761",0.00139698098425223,0.00819262048735303,0.00889328392639532,-0.00208323836270718,-0.00548816813112218,0.000673142509234337,0.00478274422141012,0.00419342095330921,0.0132889912914882,-0.00315212641401641
"762",-0.00932639701825855,-0.0137893721256525,0.00685606466815258,-0.0160056792862069,0.0171174710720616,0.00719030195922032,-0.0168760619131056,-0.0105787483516736,-0.0209127163653118,-0.0213438275954736
"763",0.00844603762114682,0.0114854648359826,0.00583620355883974,0.00306489726027892,-0.0116246000673866,-0.00479589256640345,0.0187064691149446,0.00815974177082168,0.00950314977831757,0.000807826564948932
"764",0.00270451040690611,0.000493450093608461,0.0145072092162484,-0.00258531155303754,0.0140019725934777,0.00470650007636442,-0.00345653465612616,-0.000279096524820943,0.00439302488440885,-0.0052461774260445
"765",-0.0112239524289328,-0.0180115430041637,-0.00190668163147556,-0.0115455402537873,0.00618634693827369,0.00446207251590924,-0.00910463689046437,-0.0117252265674295,-0.0104436134110829,-0.0113589960663488
"766",0.0124955289359894,0.0105532137200011,-0.000955063082183738,0.0202617360636141,-0.00285476648786454,-0.00177676725489961,0.0199082664915196,0.0155367663850481,0.00595341867261934,0.00656544367339817
"767",-0.0101686305271488,-0.0256091844262306,-0.021988581926255,-0.0240651438769425,0.01013045270066,0.00344840387625744,-0.0102966160432497,-0.0255912684617307,-0.0231348194889208,-0.0187525843160991
"768",-0.0192289896133714,-0.0308753244324098,0.00488763558224159,-0.0301650567713664,0.00457755072875243,0.00365872623848018,-0.0283915136029165,-0.019126160959933,-0.0144115932731488,-0.0124636054323451
"769",-0.0222916841402255,-0.0234331747182545,-0.0107007284351669,-0.0222169717116112,-0.00173527710254651,0.000883466501685914,-0.0229756842290617,-0.0189174471508874,-0.00186276422102727,-0.010517487817516
"770",0.00512739532172435,0.0175246766418575,0.00786655989406615,0.00732145959738428,-0.0045655064325999,-0.00220666158113259,0.00730600544665205,0.0201722166439404,0.00289264725002591,0.00467680669095438
"771",-0.00419073134485304,-0.00370948387688552,-0.0107314708608913,-0.0208022068321158,0.000327515006151469,0.0019904096285992,-0.00861291301201694,-0.0136672670453735,0.000744277984435771,-0.0110028558895792
"772",0.00475744956800184,0.00505330304781038,-0.00591736491230221,-0.00255921939922499,-0.000545762965124319,-0.00231797732271832,0.00914513604213996,-0.00353758832093853,-0.00957604145734536,-0.0145486749141351
"773",-0.0114721447815348,-0.0254038168486823,-0.00992070691609148,-0.00692824818898063,-0.000545957979599998,-0.000331863588580505,-0.0095153768306192,-0.00562131815315203,-0.000469313812722416,-0.00347368256874803
"774",-0.0108688526410335,-0.0119466522643604,-0.014027874281169,-0.0108530897738014,0.00874183672563467,0.0038737226817378,-0.0066331869823838,-0.00684311493234557,-0.00488358363400876,-0.0113289556147773
"775",0.0155508085540903,0.0200604061746383,0.0101624336550707,0.0269071741294749,-0.00907708861012424,-0.00342947304437746,0.0181904461372473,0.0161771294970137,0.0225556721645497,0.0242397840215776
"776",0.0121034047894655,0.0161636790572859,0.0191146462878404,0.00814057887846298,0.00285197084578726,0.00166611495056457,0.0165082052420646,0.0232904823634725,0.00719888338161301,0.0215144674378465
"777",-0.00498261588703397,-0.00954396392874013,-0.00987171168366763,-0.00580387984218389,-0.0115963821977084,-0.00476561621387261,-0.0115684359668694,-0.0149810556693377,-0.00394025485036897,-0.0122155473463933
"778",-0.0308661611271805,-0.0455033080882253,-0.0189429241045059,-0.0451776099517589,0.015827809575323,0.00823948176733258,-0.0373623881271643,-0.0266162969411787,-0.0398343525253271,-0.0332622435452573
"779",0.0020675012600051,-0.0190688586188542,-0.00203263108333762,-0.011164136820584,0.00217916262321616,0.00320216492595682,0.018704951270518,0.00120187263797766,0.00297017333610694,-0.0127923788437495
"780",-0.00721989560814429,-0.011149087465091,-0.00712832212329262,-0.00994629829146743,0.00130426625820013,-0.000880060100729829,-0.0227220287594471,-0.023709551319519,-0.00611386129155522,0.000446913439102747
"781",0.0125603732473902,0.0361373664837497,0.00615369664012544,0.0325818409073755,-0.00998884736097394,-0.00539946218978749,-0.00305328455067377,0.023055763247283,0.0131680410114567,0.0178651962283896
"782",-0.00195848513003738,-0.00530115278220544,0,-0.00262927099704968,-0.009541310756219,-0.00276913877881735,0.000706961608843759,-0.00120176503489466,-0.00275117151119741,0.00394900110499585
"783",0.0104664071029812,0.00729299664866079,0.00509686268319398,0.0263641467078708,-0.00542613387270297,-0.00122183758296035,0.00870957721419918,0.00721996633250011,0.0191209469428955,0.0118007183910438
"784",-0.000832622342750944,-0.00863264273103803,-0.00608516566833883,-0.0125866367909269,0.0041196573837905,0.002335270135434,0.00910172352746463,-0.0062720986670286,-0.000840063497808186,-0.00561547411050289
"785",0.0157351125576002,0.0230338859271666,0.0102042775995432,0.0257545044711018,0.00188493754705088,0.0022200751569792,0.0268269087226505,0.0135253570441207,0.0241031574728778,0.0304082808699191
"786",0.00473828780125363,-0.0010984796281841,0,0.00355074099339081,-0.0113989948014467,-0.00531563367648635,0.00945989491649546,0.00207592539837242,-0.00337532375364014,-0.00505895277612167
"787",0.00589553464395287,0.00494791886520707,0.00202007303541007,0.0037906497931508,-0.00403033092103122,-0.00356117022249058,0.0133864573895184,0.00562308774108899,0.00668194965675051,0.0088981828450192
"788",0.00207355959071021,-0.000547061944684346,-0.0161290784478111,-0.00855999227191295,0.00539503237998762,0.000558870619595808,-0.000219764040646941,-0.00971151679145565,-0.00463722482349815,0.00588001847142516
"789",0.000180050801480647,0.00136836610571844,0.0122950267949173,0.00126970945006866,-0.00413624839619853,-0.00078198461917256,0.00418377478815946,0.00267459863993214,-0.00365397822550495,-0.00542802922543661
"790",-0.0121448215841334,-0.0210442808351411,-0.00404832543598077,-0.0230789049468008,0.0156039832951356,0.00759776308894899,-0.00789482915677031,-0.00859516256301351,-0.0108187494269734,-0.0163728741687471
"791",0.0091978536164079,0.00949237483983523,0.00203227020252861,0.00960539708609764,0.00243172800167213,0.000554890877738856,0.00972618171404016,0.00956638272146959,-0.00491239229689866,0.00810937083926322
"792",-0.00135359827245995,-0.00884996575694885,0.00202838855611298,-0.00822839949529008,0.00562353431969864,0.00365688388343188,0.0050343042498362,-0.00444193101865697,0.00884870520819003,-0.0169348735900949
"793",0.000632283140601819,0.00502269800625466,0.0060729673804325,0.0101114313265369,0.00515350033633366,0.00154581468506509,-0.00239542904971601,0.00832861383520056,0.010340707420196,0.0176571726432413
"794",0.0103850380844099,0.00222078770374612,0.0100601975647618,0.0169406235355209,-0.000437465737403775,0.00103955734159866,0.010262281887969,0.00855485985442006,0,-0.010156572821003
"795",0.00277059661135559,0.0132962213499654,0.0029881084601433,0.0113580687623267,-0.00131370419557342,0.000552794983982974,0.000432193269085834,0.0152089010628293,0.0145298090103263,0.0106884025606933
"796",0.000891042100767514,0.0120286361696917,0.00695170659032285,0.00124759752343673,-0.00252197388844932,-0.000993908684689293,-0.00216080429148158,-0.00316938195452754,0.00549450564297893,0.00972926960187404
"797",0.00302786767064656,0.0013507714474652,-0.00986235267690994,-0.00523417125091563,0.00527573863731212,0.00176762507515238,0.00411380329405153,-0.00115591752719657,-0.00716648769595518,-0.00879774891871954
"798",0.0142932300992125,0.0207711977869469,0.00996058750374096,0.0260583939135171,-0.0131190162514043,-0.0047424813662178,0.0228545518047181,0.0205438835302951,-0.000180492643138241,0.0118343758967849
"799",0.000174976116454229,-0.00396417588430453,0.00690313032318923,0.000732890165198619,-0.00520663756185691,-0.00265967369342812,0.0124370980207082,-0.00481992348757276,-0.00839275351308999,-0.00125311570013642
"800",0.00166269786698758,-0.00159158285368544,-0.00391802865316215,0.00561219950328451,0.00022262606957546,0.002556320471514,0.00333091060504387,-0.00113924731221204,-0.00145609760073084,-0.0108741776279682
"801",0.00445569682072944,0.00425197826686063,-0.00688279980640794,0.00703741100985433,-0.00256059846114365,-0.0016635639796293,0.00539577153422122,-0.00912753975660319,-0.011392635696385,0.00295987758725458
"802",0.00417514345936931,0.00846762589434302,0.00990082880813858,0.000240611033167193,0.00368350904077674,-0.000887715150863833,0.00495339100526571,0.00690843091015014,0.00119846039274951,-0.00252956316850506
"803",0.0000862996865320653,0.00472338013349272,0.00980387947278727,-0.00337249131827644,0.00622774105799428,0.00155577116492567,0.00739328042349552,0.000571808114484984,-0.00598527635332002,-0.00591707919774553
"804",0.000260003389239927,-0.010707854950989,-0.00485407535270144,-0.00725164975668546,-0.0013266493866434,0,-0.00285415978270986,0.00171459748320046,0.00379809181467605,-0.0119047301272583
"805",0.00796616189567012,0.0163673425615123,0.00975616868091134,0.0129047638231108,0.00796811539342168,0.0038827185481094,0.0259658680568464,0.0168280811140986,0.0188261441599655,0.0133390202979642
"806",0.00592736818311712,0.0028573686588107,0.0038649451861863,0.0108174693630609,0.00428231634265086,0.00121629442589066,0.0121563619217278,-0.00112207290324784,-0.00733701073664839,0.00891716287918798
"807",-0.000512395878424665,-0.00699314025266029,-0.00673728603206947,-0.00760986877354575,-0.00328061730618812,-0.00264962415683401,-0.00393757260319727,-0.00224671701160439,0.00684369036750399,-0.00210443502469138
"808",-0.00506162339895166,-0.0112153421819391,-0.00193852003383477,-0.0129407461844578,0.000987688783145702,-0.00132807758698938,-0.00849975194166264,-0.016198899314217,-0.0186695402816581,-0.01223100333295
"809",0.00534582099129577,0.00131887971559896,0.00485473615027887,0.00364204650849298,0.00109634912953527,0.00332443740863875,0.0103666146173809,0.00660946455038824,-0.00489470820922344,0
"810",0.00703332432540904,0.00579559988511491,0.00966190550106361,0.00701479892362755,-0.0047069557176953,-0.00209934819560798,-0.00276201039240553,-0.002569381205621,0.00529002320185601,-0.00426988417232754
"811",-0.00485483340667892,-0.0154531034148161,-0.0162680220906961,-0.0148931234035464,-0.0182555191013555,-0.00996054659946632,0.00316580966778357,-0.0151683545109769,-0.0186484213441653,-0.0111492962624892
"812",-0.00162599307973232,0.000531890362387655,-0.0058365489934179,-0.00268224412773288,-0.00638552452529306,-0.00368890778862596,0.00157358040243016,-0.000872496197010575,0.00451548435045668,-0.0056373907344931
"813",-0.000600064131510258,0.00771079646157746,0.0156553889488664,0.00489011905720727,0.00281855932126907,0.00235642787774215,-0.00357965919715098,0.0116348343811705,0.0169507119025165,0.0017444157174622
"814",0.00634751023045665,0.00949856269071181,0.0125241858778848,0.0180047074997558,-0.00382342734844077,-0.00145551217062212,0.00439049734884156,0.0212767931259361,0.00147346906615597,0.0226382280421098
"815",0.000681854631978673,-0.00444309232632623,0.00570893538107065,0.00382409149501983,0.00316158596925709,0.00100877149842526,-0.00198683976322944,-0.00281557961077317,-0.00717240459770119,0.0021286238789695
"816",-0.00340717081681208,0.00656330746946332,-0.0122989723237916,0.00285712051530562,0.00686183271038043,0.00235173386864918,-0.00895922364152568,-0.0095989332963996,0.00907655821916675,-0.000849649729898538
"817",0.006837480453461,0.0164320147273509,0.0153258264501404,0.0261160824625786,-0.0024447141919165,-0.00207202508786897,0.00462061323052776,0.0193841349213275,0.0120239103815671,0.0195577740490089
"818",0.0081497442489451,0.00538853270081163,-0.00283032871293554,0.00902331996890338,-0.0166382799654207,-0.0089832136183795,0.020795724699689,0.00531316571907681,0.00571374014667625,0.0158465370998924
"819",0.00235753835723052,-0.0068911255331997,0.00283836221099909,0.00298115063985716,0.0015995837896241,0.00294585693460392,0.0201767277990985,-0.000556251682812592,0.00126251241106057,-0.000821006858102935
"820",-0.00571261780878229,-0.0110513270633112,0,-0.00868767374554125,0.0127840867800117,0.00621376530239504,-0.0215057089022928,-0.0158641792045926,0.0131495903192793,-0.00369756658899045
"821",0.00346423444615596,-0.00051944657495695,0.000943238178234607,0.00345920346484552,0.000451489683787498,-0.00112268882271171,0.000392276198765362,0.00735308833793646,0.00142238423721897,-0.00164954680753537
"822",0.00656722900876261,0.0145605458233964,0.0028273268639869,0.0062056712084344,0.00236549230886807,0.00112395066956572,0.0158891803477341,0.0106678446594868,0.00878825550309359,0.00206531912904606
"823",0.00158937188260566,0.00794473591017342,-0.00187946843781006,-0.0079944474872774,0.00528230763428161,0.0026939196920519,-0.00656543227574735,-0.000555231578312054,-0.0055437962473055,-0.000824475860280893
"824",0.000751795847694137,0.000508254819752585,-0.00188311894944149,-0.00207243346733488,0.00324240031263567,0.00190350285370933,0.0227406469852671,0.000555540031680568,-0.00283160777220404,0.00371290560147886
"825",0.0113492008177094,0.0142309476027704,0.0047169167381742,0.0147669283806418,-0.00702123911571773,-0.00268211693173537,0.000950186750848792,0.0127779518842543,0.00301709995532695,0.011508480076293
"826",0.000825215532389789,-0.00350755226270305,0.00469485524844671,-0.00545695491438591,0.00112252665757673,0.00168134605525139,-0.0248715515156672,0.000548421936290566,0.00548529598766079,0.00365708345691451
"827",-0.0159122917214691,-0.0213730408334791,-0.0186916110134629,-0.0292636849831265,0.00728656804779271,0.00603974569118781,-0.0208332633940718,-0.0216555570741785,-0.0212054901679632,-0.0182186646443475
"828",0.00376992310256608,-0.00385417329035109,-0.00190495022136672,-0.00400406430916056,-0.00244931615708388,-0.00244551156086159,0.00377763376726481,-0.0050434842371202,-0.000809025544930342,-0.0127835421184697
"829",0.00893078517396861,0.00851195270653071,-0.0038166919386583,0.0118235176739541,0.0035709969964679,0.000445576769492417,0.0156499980776252,0.00816654326659028,0.0027889968009176,0.00793648541716063
"830",-0.00181967097022173,-0.00818413941884422,0.00383131488730304,-0.00327183818394616,0.00822556543740616,0.00323156074058306,0.0187241711782313,0.00139675479451995,0.00762604528643496,0.0049731226595251
"831",0.00298338489140804,-0.0108302208357638,-0.00858747921061043,0.00422023358392698,-0.00297711592139527,-0.00233231574306392,0.0145512034487201,-0.00223141209262667,-0.00418486339924962,0.00247419288560891
"832",0.00652767251339248,0.00860235815517729,0.00673702969905632,0.00537001778219226,-0.00353811769631962,-0.00278317671461259,0.0130210626969032,0.00698918118647152,0.0120708695304317,0.00658156363703033
"833",-0.00377647862193464,-0.00155037561759419,0.0066919741518956,0,0.00110904754240626,0.00066996368921135,0.00633405597751202,-0.00111044014664263,-0.0038872867941111,-0.00490381329421719
"834",-0.0236502957170267,-0.04452522165489,-0.0180438718220668,-0.0357640985954766,0.0140782765092138,0.0093710170320096,-0.0316549731613667,-0.0330740284713151,0.0166740310421287,-0.0151951590075315
"835",0.00759638976383625,-0.0048768339348676,-0.00386845556812465,0.00842968835653268,-0.00852602847192507,-0.00508457928303618,0.00344123122441986,0.0063235538482278,-0.00279158168345772,0.00333606789495611
"836",0.012397275083879,0.0185137270872373,0.0116508668529367,0.016479339022041,0.00418952824337238,0.00166646178002194,0.0413412338063597,0.0159956724636672,-0.000262435487051516,0.00789703081839277
"837",-0.016961877985084,-0.0155039659178241,-0.00287888077081111,-0.0119827801643418,0.0115283846860545,0.00609985561167803,-0.0311015600589999,-0.00590403991908561,0.00945049010719701,0.00783502902155764
"838",0.0129618439538943,0.00705978133242868,0.00288719265422488,0.00546962818016938,-0.00130733356791402,-0.00262048082623212,0.0309662512422302,0.0152717600764867,0.00320736821075451,0.00490995854541798
"839",-0.0235146176559602,-0.0401728026472596,-0.0307103429779005,-0.0458845542879978,0.0179959477457299,0.00676212040273394,-0.0234426897453909,-0.0406686241204169,-0.0074310894124836,-0.0268729322961048
"840",-0.0059564710122415,-0.0269663172952976,-0.000990050651648811,-0.0180963234719201,0.00589213644987119,0.00385336798377844,-0.0140657406342565,-0.015389186958487,0.0019151475080923,-0.0225941773588147
"841",-0.0332135486528448,-0.0534062238168374,-0.00594654287943741,-0.0408985234836415,0.0308868271549481,0.0109682681705552,-0.0401372207115298,-0.055145896708145,0.0295421158933744,-0.0196918202787819
"842",-0.0148751684413578,-0.0057946600123373,-0.00897299665888041,0.00526407699863385,-0.0125010481260495,-0.00271210679999545,-0.0168451547363881,0.00530574845609255,-0.00185670523852988,-0.00524014825566066
"843",0.0440409831184339,0.0763806420543554,0.0281691247817759,0.0720087033534449,-0.0207158228646833,-0.00761514374551331,0.0659138282119109,0.0509158824216644,-0.0059186354760794,0.0193151962987981
"844",-0.00284093636960236,-0.00541480560360064,-0.0225050631809997,-0.0180752262793759,-0.00256370009569507,0.00120621080291627,0.00113485232024235,-0.014180149854548,0.0262822488730119,-0.00172262936785217
"845",0.0139859336859156,0.0163323084702338,0.0090091317662464,0.0124378827270279,-0.00760486675607086,-0.00251918846018706,0.0162451611125269,0.0107881425304912,0.00613291874248567,0.00819678682120339
"846",-0.0124304364748025,-0.0219902511337501,-0.00793658901876981,-0.00933694635818849,0.00658321344104618,0.00274459807742722,-0.0131973269085525,-0.0103765166926297,-0.00691930795849582,-0.00855803888595574
"847",-0.0181051429535234,-0.0302683811017076,-0.00699980575658876,-0.0205850305379569,0.017371245310728,0.00645866535474693,-0.0308909835294038,-0.0170756098313831,-0.00157593731877792,-0.0254639689982534
"848",0.000526583878657449,-0.000594385523936869,-0.00201429784322427,-0.00607765973522578,-0.00368911411784134,-0.00217498107675085,-0.00155470525118229,-0.000305286293781126,-0.00839081145491039,-0.0283436440301731
"849",-0.0136022360440495,-0.0190364805481604,-0.0171545960917111,-0.0208914796826583,0.0153393531828814,0.00730309790089789,-0.0255011640219898,-0.0216464026873832,0.00108911694797986,-0.00136734681240436
"850",-0.00569399179720065,0.0042451222422113,0.00718699463049721,-0.00962805206696382,0.00333429727433932,0.00086546331571391,-0.00839031652996425,-0.00218156446925188,-0.0239350660964945,-0.00912836160459607
"851",-0.0377593864849172,-0.031400858566577,-0.0152902863958163,-0.0496584456700644,0.0210796016858814,0.00973096757115566,-0.0483477832030885,-0.0371640053426897,-0.006773566152111,-0.0207277302351985
"852",0.0145990180002686,0.019950325771708,0.00931668085367865,0.0323472113794752,0.00101713005601822,0.00053547788339614,0.0323875166813905,0.0204347748155094,-0.00535216696658036,0.010348075457902
"853",-0.0128311827427818,-0.0259782498730183,-0.0133332269024754,-0.0104443746555223,-0.00345470938364245,0,-0.0200942202975313,-0.0171647227264558,0.0140600155002604,-0.000931085981564328
"854",0.00102139289169423,-0.00156887674738249,-0.00623731544732375,-0.0108254879844778,0.00489299560690504,0.00342449814642398,0.0104625339763846,-0.00840884846886669,0.00445057358612022,-0.00792165449983961
"855",-0.00602866891979559,-0.0141421208024761,-0.0125523702870302,-0.000547343890177965,-0.00283922853109186,-0.00202664147604104,-0.00393421314958819,-0.00913220823504579,0.00945807762902118,0.0108030940099144
"856",0.0334981794511489,0.062161432063881,0.02436459994664,0.0604983373916368,-0.0226886313066186,-0.00951102398561698,0.0542615905904238,0.0513495266596544,0.00185701863883669,0.0292750765132741
"857",-0.0125493597821262,-0.0204083104143357,-0.0165458220266219,-0.0165201666371122,0.00458048863663385,0.0045313395611426,-0.0149869282962247,-0.0159677474985794,0.00160076667620235,-0.00857780778638462
"858",-0.0168238872082817,-0.0119483793477242,-0.00315485497039547,-0.0183728639206073,0.00702892390420851,0.00129256901092378,-0.0194195122932732,-0.0104993819589173,0.00866425829401729,-0.0186703822178462
"859",0.0260392775698954,0.0310077289699191,0.0052742852125196,0.0350268167889016,-0.00949880918615009,-0.00570136442095937,0.0220497814220539,0.0369773260881303,-0.00108418810493904,0.012065039772875
"860",0.00344419338840085,-0.00210528381447672,-0.00209837818720082,-0.00361687974543179,-0.007297248415577,-0.00140634133909745,-0.0025970048381907,-0.00279081105147905,-0.015194523419557,0.00550208235748162
"861",-0.0351370438872997,-0.0491259806092536,-0.0189274183897111,-0.0355195667548482,0.0268818381048264,0.0138676903288582,-0.0542758426787546,-0.0407334394802956,0.0104272889998924,-0.0310077024594181
"862",-0.0124504552993839,-0.00919176915077369,-0.01607745944303,-0.0155913892698063,0.00766996515021123,0.00406067586518266,-0.00508255290293502,-0.00842810117465742,0.0192968869989614,0.00188232704909397
"863",0.0107118162804809,0.0111963526931662,0.0098038943896348,0.0229381007174767,-0.00497312571051323,-0.0030868601618933,0.017453941019473,0.0117686212135992,-0.00403323736987793,0.00798490818368358
"864",-0.00534606413494843,-0.00284706806487323,0.00107904718110019,-0.00533892017657112,-0.00112148809712409,0.000107225943740019,0.00502088301589532,0.00387720552529869,-0.00363638016528933,0.0046598644724829
"865",0.0292312814124942,0.0491751807077392,0.0172409796085644,0.0348898341633403,-0.0178682010094799,-0.00928655193845274,0.0418402710407766,0.0379786321677353,-0.0131884292167954,0.0166975025710112
"866",0.00485621619705445,0.00332616841463773,-0.00211838418731236,0.00518655275369939,0.0126836690316781,0.00635691076520351,0.010389831181695,0.00186054070098596,0.00874170792013351,0.00136868840960847
"867",-0.00155009063194123,0.00693192545096677,0.0063692720813957,0.000258163823395385,-0.00513358936570596,-0.000856414143217576,0.0118640813852735,0.00185736137720061,-0.00341641524178959,0.00273344776777806
"868",0.0227374008103509,0.0359173390445258,0.0179324573469917,0.0301778719282351,-0.00412725433025563,-0.00310762040465207,0.0216927436870795,0.0299653502095947,0.0116220737729444,0.0168104514110876
"869",-0.000356785409180937,-0.00953474134930143,0.00414542759324199,0,0.00569860360727747,0.00279484547978925,-0.00726853021658525,-0.00419895742795162,-0.00545496331027306,0.00223419928982249
"870",0.00160707164863405,0.0055424739096126,-0.00206421806117041,-0.00500765867900732,0.00813901644744397,0.0047160157709123,0.00154167929038751,0.000301485526305267,0.0130474526211677,0.000445917171275401
"871",0.00108462189694913,0.0011603446541617,0.0020684878711934,0.00452964086960139,-0.00163456906028914,-0.00202643261545843,-0.00288599707674997,-0.00671323728568096,0.00762920414062007,-0.00178259847966811
"872",-0.00286405211025165,-0.0066301228960669,0.00722370962092733,0.0172847837120962,-0.00286587390745818,-0.000749164504219912,-0.00713866350091563,0.00214055776306821,-0.0198648779636101,-0.00401780231396276
"873",-0.0165154854431121,-0.0092371232344719,-0.0122950267949175,-0.0192073196039388,0.0119076885949443,0.00599178113950294,-0.0281772789647325,-0.00762879719008247,0.00880470146029322,-0.00224111676075323
"874",-0.00310323607516472,0.00661631235987414,-0.00428390516021582,0.0025779697300532,0.0067974941644342,0.0037219206261796,0.000599606648844508,0.00492008749816897,-0.0041169206451277,-0.0166218384377776
"875",-0.0165703759615716,-0.0179264330753711,-0.00314755893541763,-0.0176454858599372,-0.00594488929975823,-0.000847717237204337,-0.0205997014541995,-0.0140758950371839,0.00289380743018963,0.00228421090344666
"876",0.00418908302651055,0.00212945971876044,0.00421033665343318,0.0118038208693199,0.00405445529183801,0.0015909635234026,0.0255195631692104,0.0117938780119384,0.0120362651598616,0.0182315253844831
"877",-0.00315222221927502,-0.00394629581263028,-0.0115305817495008,-0.0068474683239369,0.00938941213390487,0.00709392081425553,-0.0114384528055114,-0.00797532577350879,-0.0136038283870344,-0.0107431451285394
"878",-0.0308749009663637,-0.0374887643472092,-0.0243900812815773,-0.0406027975237921,0.0109019349955148,0.00430911862804351,-0.0320747778134657,-0.0281385420944603,0.00148650595380317,-0.0276017606022768
"879",-0.00949995528065894,-0.00728318059470523,0,-0.00665427745509228,0.00672831470421875,0.00146593427218478,-0.00985737870065007,-0.00827226712789064,0.00338091044893818,0.00372261089084946
"880",-0.00445656624986612,0.0169061060746849,0.003260779244038,0.00723457833911234,0.00157706984153427,-0.000439818085931409,-0.00190650868627729,0.0134742780326778,-0.0381327991452992,-0.0152989615223466
"881",-0.0054497741779409,-0.00470505248845987,0.00433359604882688,0.00425668599686779,-0.00797250686566242,-0.00178275331765754,-0.0190999846823321,-0.00158271828705281,0.0123889011244966,-0.00188311652441298
"882",0.0065559502369994,0.0226914860516043,0.0204964423065161,0.0185429520139306,0.00823534877705345,0.00241591848683242,-0.0194718660175792,0.0117310962882409,-0.0167102374328676,0.00283005256186408
"883",0.0314961098951763,0.035439031738546,0.0190273293157737,0.022106361460281,-0.0117101479747119,-0.00314312483292323,0.0476607433289793,0.0363522880365899,0.0104712125916879,0.0225775443640059
"884",0.00989545568789585,0.0104166090807618,0.00207485509570193,0.00483493360060661,-0.00637316450507908,-0.00241730808270635,0.0107412934799795,0.000302387870286802,-0.00441691995879756,0.00919974372801868
"885",0.00746555337332455,0.00147279097688524,-0.00621103825281544,0.0121550516559297,-0.00571202969421958,-0.00263395661997767,0.0131274947067044,0.00030240329691722,0.00981146668212163,0.00182312908320581
"886",0.000647990502615325,-0.00264706221058009,-0.00520856557758476,-0.00800598190028512,-0.000402699948474639,0.00168999070142806,0.00370234941406045,0.000906401604853446,-0.00861781844695997,-0.0113739613018505
"887",0.0150886550557832,0.025361278527138,0.00523583677679018,0.0116011367164575,-0.00857062834267308,-0.00495695808592544,0.0219263781833996,0.0132850349800788,0.00869273082300093,0.0161067811886209
"888",-0.0000913317880164577,0.00258832625885907,0.00729123893555883,-0.00199430295626224,0.0100683423235586,0.00498165192571998,-0.00581503988307219,0.00327754306955175,-0.000506911114338315,-0.00181156937638549
"889",0.000274020390821805,0.0100401445545906,-0.00827288343892318,-0.00474636110008908,0.0099679812757989,0.00516747037360177,-0.0022190694395281,0.002079363129176,-0.0005917159613259,0.00952804655642714
"890",-0.027534628786004,-0.031241037165498,-0.0250262057116579,-0.0298696724612302,0.00488463670222505,0.00577110052312202,-0.0307255656456462,-0.0222290471050116,-0.013194662610302,-0.0125843292251807
"891",0.00590621818793879,0.00586353004818196,0.00320859379001504,0.0131956543954381,-0.00615091781461707,-0.00260785312377865,0.0114704510544126,0.0142467499772352,-0.00805686994183386,-0.000910226211123244
"892",0.0110916485913066,0.0020400853658431,0.00639647535145316,0.0234932891497703,0.00149707998766768,0.00104595599361357,0.0171134050743709,0.0140468423836104,0.00794952887022737,0.00820039019244789
"893",-0.0129982310251837,-0.0171611967605598,-0.0180083344553296,-0.0102295439225429,0.0169445789288849,0.00637279574306948,-0.0192582504386762,-0.0132625024920511,-0.00685815676196899,-0.00271126125667331
"894",0.022322149018819,0.0361052424181281,0.0183385817692669,0.0302493732955955,-0.0115657624963567,-0.00550201384012838,0.035965336218106,0.028076365755644,0.00871819609353808,0.0199366670670988
"895",0.00867916926343892,0.0131392663680592,0.0148308910542014,0.00685069811220451,-0.0106095623002957,-0.00323632227585191,0.011771699826377,0.0136545488671933,-0.00658912368142117,-0.00310973207646137
"896",0.0104155470478364,0.00733019364271992,0.00104367947818407,0.00680465384803197,-0.00170375792482802,-0.000314247501316589,0.0258335972296888,0.00917175538960269,-0.00490997518855973,-0.000891345105075714
"897",-0.0000896001817540792,0.00643724623674902,-0.0052136307383539,-0.00168922011123784,-0.00963742781206745,-0.00345715348435549,-0.000192421891696104,0.00198816565909188,-0.0173995416568441,-0.0107046737841719
"898",-0.00645459830477546,-0.00834292221567023,0.0115303353728393,-0.00556108951357615,0.00324337142756193,0.00431035895113063,-0.0015384353479877,-0.00935341051800742,0.00237861858199961,0.00405774690872085
"899",-0.00487221805279581,0.00224349657492784,0.00621744463123086,0.00170187009942291,-0.000302164308552455,0.00209324005347788,-0.00885797323661675,0.00457774985039117,0.0044823519465842,0.0143690478374703
"900",-0.000181453143848098,-0.00167885592368122,-0.0082387731001311,0.00485440403752935,0.0155648711162313,0.00585013145997726,0.0034972286508923,0.00113952436823617,0.0104995799238814,0.0132802587701601
"901",0.0225808344401661,0.0369957069071432,0.0218068915052818,0.0258455044417902,-0.0140383090636388,-0.00309233694412248,0.030396986411088,0.0301560111961632,0.000432963900475647,0.0192223290506586
"902",-0.00478866232248631,0.00135109623930485,-0.00406530633937752,-0.00470921096966548,0.00577186824296305,0.00470010144737487,-0.00526111406158858,-0.00856099738698901,0.00389472906443888,0.00342901439923127
"903",0.00668329176839033,0.000809765926394368,-0.00204059049739302,0.00141931669959838,-0.00765159370319501,-0.00415859908123029,0.00321104146973328,0.00334275486395419,0.00629367197678543,0.00854337299574337
"904",-0.00106235838147428,-0.0002693191631018,-0.00102257677932682,-0.00448835094113409,0.00466645837128277,0.00480147016013333,-0.0124267694083161,-0.000278015044209878,0.00222757023451359,-0.00465902280095076
"905",-0.00407651791684271,0.000539468355647887,0.00921179967051233,-0.00142392887093001,0.0109069615154469,0.00654576293091269,-0.00324115075894404,-0.000555301415900877,0.0073516240207312,-0.00893604810459558
"906",0.00533893315279599,0.000808640127364812,0.00101448875038157,0.00522821522860339,-0.00369629138396377,-0.000206252710011845,0.00994645102235592,0.00611278960481076,-0.00373382565287939,0.00343490326253937
"907",-0.00539880742128818,-0.00673475897899767,-0.00607909666207229,-0.0137117565791233,0.00210631559656194,0.00505892782944772,-0.00776547334097577,-0.0107703736179992,0.00281091136608325,-0.0106975486074448
"908",-0.0274068894235021,-0.0461080105994043,-0.0336392001494358,-0.0318789564654891,0.0134071374692577,0.00564969968656936,-0.0240502871313318,-0.0337799488471114,-0.00331272394514415,-0.0224913537169457
"909",-0.00612991323372281,-0.00255907840196878,-0.00316465543028854,0.00173283699742788,-0.00246813661448053,-0.00255346585163674,-0.0115392791299602,-0.00115562932757884,0.0121868165054311,-0.00752215774694576
"910",-0.00294603289210693,-0.00427574333243375,-0.00105837917819129,0.00543730778103391,0.012472058654718,0.00430076097356746,-0.00217660090570715,0.000867494740516062,-0.00025258062438116,-0.000891650799776267
"911",-0.000461829398832325,0.00601181420845931,0.00741585013044088,0.00934137793912337,0.0250262120921687,0.00723983194688627,0.000991603845195588,0.00289031747476343,0.00833758646349314,-0.00312356292659821
"912",0.012285433366787,0.0108140753080876,0.00525727059329606,0.0104725582266729,-0.00572219303479482,-0.00506154740094156,0.0217907795496304,0.019308140661447,0.000167017451757623,0.0143241167204717
"913",0.00182511361942961,-0.000844758617768115,0.00627646907709245,-0.000722895906580256,0.002685964822702,-0.00101789275167852,0.000193978409364526,0.00452359356503029,0.00392485177453028,-0.0039717927589521
"914",-0.0173970525835336,-0.0166243064215872,-0.00207904582687468,-0.00771858617210119,0.0155937145847531,0.00448201516591418,-0.0226788660558476,-0.0115393095234081,0.00141405754937574,-0.0101905157808873
"915",-0.00324433715649741,-0.0160459631267127,-0.00937492224519831,-0.00291672295393508,-0.00113109677935652,-0.00324492003203425,-0.00297502437120611,-0.00740341606021866,-0.00348864526529324,-0.00626679242697858
"916",-0.00381268080033792,0,-0.00630955885608198,-0.00902005184312504,0.000189275636480302,0.00132211621811518,-0.00477438780390649,0.0014344056102864,-0.00158374592328292,-0.00675680343109109
"917",-0.0148433816052592,-0.0171811490289855,-0.00105837917819129,-0.0127918689910149,0.0160287316964263,0.00792444883889631,-0.0043973156145225,-0.00887999938447925,0.00484222745735696,-0.0113379006567939
"918",0.00388538077831257,-0.000888863724192057,-0.0031773500311264,-0.00647905603152288,-0.00324803389996109,-0.00453552731660678,0.0130496340813155,0.00780339242669714,0.00830840803997668,0.00504599179799725
"919",-0.00670175569029385,0.000296670392021525,-0.0010630025560332,-0.00627037677134445,0.00940311147634487,0.00455619205010982,-0.00554890957595822,-0.00286727903530504,-0.00329599535847069,0.0114102993379197
"920",0.0154896908861659,0.0195671885727267,0.0127660728936296,0.0219585725128628,-0.0283159657940016,-0.0114906736100855,0.0159426654992085,0.0192693140121976,0.000413384593364707,0.0171480117157852
"921",-0.0145049537974422,-0.0171562053983775,-0.00315145066722855,-0.0165470452892893,0.0191742748163872,0.00764790595698561,-0.00921949928009802,-0.00846533119361137,-0.000826361444072998,-0.0017746899064317
"922",0,0.0056213001258556,-0.0115912723495912,0.00602681705408292,0.0110833939380093,0.00445213149004253,0.00930528938892028,0.0082527280286806,0.00967660211143473,-0.0133332888102071
"923",0.0299117689774591,0.0385407525877279,0.0277186445413491,0.0351972316667364,-0.0206768634853556,-0.00720017289223285,0.0315806017853482,0.0273782412879864,-0.00319462642210622,0.0198197805590823
"924",0.00931220284687306,0.00821525317044869,-0.00311188643455351,0.00168791689133529,-0.0105661123199284,-0.00417138961294872,0.0125504804112666,0.00576906524452769,0.0049305529635868,0.00706713234755285
"925",0.0129715776436417,0.00983405658438685,0.00728374469279913,0.0117956565944448,-0.0123947210068448,-0.00572101978418538,0.0131449613652059,0.0106530817393677,-0.00351623187900707,0.00526322156738601
"926",-0.0112723665374115,-0.0178072517813107,0,-0.0145131016886718,0.0204667281603796,0.00791157092333372,-0.0139014278245863,-0.0132434829944293,0.00689312319962965,0.00523562019718837
"927",0.00702307791385959,0.00736534326256466,0.00206637275111121,0.0108641107794851,-0.00794612801467043,-0.00275241648132196,0.000563857624343411,0.00520408495646185,0.0000815158944136307,0.00217010912772109
"928",0.00461906163070114,0.00899877047618625,0.00309287974327921,0.00573206330402098,-0.0197412083221969,-0.00787075956479855,-0.00751428578094582,0.00844679027217965,-0.00937169757453915,-0.00563024417114466
"929",0.00504876406695387,0.00641044788404455,0.00719391418949722,0.00356211029642384,-0.00457245999848988,-0.00288497146957278,0.00397470101243025,0.001621130454043,0.00139852749915326,0.0104531334813114
"930",0.0111226896502026,0.0160619832497966,0.0102044215082584,0.0238997735530324,0.00488597978528849,0.00475323165978536,0.0156487924878963,0.014836890873192,-0.000903639179241633,0.00732757416011309
"931",-0.000620703305127535,0.00953947758999463,0.00303051571681623,-0.000462285569790222,0.00962962234192744,0.00503915975587232,-0.00297019979280322,0.000531583390435575,0.0197335466271942,0.00299525195401307
"932",0.00381720646249817,0.000539833199730833,-0.00201434811394785,0.00138727039569009,-0.0148346983639854,-0.00347951613179043,0.00781975659627054,0.00106297749658513,-0.000645016948355503,-0.00170654908078371
"933",-0.000265708586746349,-0.00215852833238805,-0.0131181338839815,-0.00507981979012728,-0.00987608053588085,-0.00349071276335078,-0.00535772390530753,-0.00371557966452207,0.00556716950835612,-0.00512813520556832
"934",0.000373511680435534,-0.0102759657979016,-0.00306745996602453,-0.00162425875175931,0.00404871860006373,0.00226674176391106,0.00297229006010102,-0.00583069285720239,-0.000722105449460941,0.00343637901994409
"935",0.0152903123752792,0.0193990146833589,0.0174359072950465,0.015806559044736,0.00580312485582812,0.00308423531953772,0.0224071503223187,0.0172969416989281,0.00264976712180998,0.00813358273024756
"936",-0.00201342324227471,0.0026802061772,-0.0110886792539446,-0.00297510595957118,0.0138862680936287,0.0093263921575788,-0.0157581446504097,0.00239139080692219,0.00912948644679701,-0.0106157845556669
"937",-0.00491322604603384,0.000267407778430151,-0.00305816900340816,0.000688696379305576,0.00896977358822459,0.00152344926645798,-0.010305490808071,0,0.00150777713661165,0.00600867863313748
"938",-0.0081114233121391,-0.0117584399845383,-0.00409003674535136,-0.00642194070641522,0.00286781416441806,0.00141990794462354,-0.0224323148043503,-0.0108666172782984,0.000792440589360677,0.000853142814789987
"939",0.0206218321336766,0.0316388706620863,0.0133472175429228,0.0184672395779732,-0.0134398061856683,-0.00496158072290154,0.0272447743773667,0.0262590473635027,0.00308787799474564,0.0153453669436308
"940",-0.00479004246466053,-0.00655327772123071,0.00506575512563967,-0.00181329425979071,0.0173909355104565,0.00773302613043203,-0.00989887695043556,-0.00626599139892181,0.000236790587468727,-0.00671712532960733
"941",0.0035007619526124,0.00897114441838087,0.00403252163510937,0.00726610147046092,0.00683793778442254,0.00333173949468923,0.00264130864636281,0.010509522256573,0.00891727423518573,0
"942",-0.00174422675260943,-0.0047072579808155,0.00501994991819932,0.00338162958681787,-0.00414980708663393,-0.00241532626057495,-0.00733819163181049,0.000519917665885883,0.000782158792055565,0.0131023214391592
"943",-0.00297061936160448,-0.00551772775132198,-0.0119879134669605,0.00584118163195102,-0.000664060183534487,-0.0012097065586294,0.00227457753629645,0.000260142436406596,-0.000312567416472787,0.00584064025226727
"944",0.00420587149678231,0.0105682267488261,0.0020220496274066,0.0147419069031023,-0.00483236817078714,0.000536494240525709,0.00491669729267863,0.0161078411863416,0.00781799678467676,0.00207379995796053
"945",-0.00750348926323841,-0.0138564080559429,-0.0191728122929326,-0.0030814915974916,0.00258079427025093,0.00354137136034582,0.00846817306579473,-0.00946023300048382,-0.0034907841597771,-0.00331121313906824
"946",0.0201315832566908,0.0291624146308411,0.0318931766441823,0.0181055196195754,-0.00600665956981261,0.000201342609894795,0.0130620714898046,0.0216829160069583,0.0196948300026172,0.0203488153415423
"947",-0.0000859243702807655,0.00566719264788884,0.0109672743131177,-0.000433705788603911,0.0125662250555374,0.00645179548170383,-0.00294692721593492,0.00757971935204638,0.00625996617070146,0.000406994849060593
"948",-0.00120648687788538,-0.00179291326378594,0.00394436415697164,-0.00889572127867255,-0.00833637752576111,0.00100171726270415,0.00221682160432923,0.000752327047804702,-0.0109248389488635,-0.0101708574073451
"949",0.00560862650671434,0.00487533727440947,0.0049119282743546,0.0120404885959122,-0.00439500146706517,0.000399891085920201,0.00129002750479823,0.0065142857945526,0.00989498388797205,0.0332921999423756
"950",0.000944047407607451,-0.00229843715555345,-0.00195496088340674,-0.000649469126167923,0.000192625839370519,0.000999839724998841,-0.00147209008553484,-0.00174268460827753,0.00478496871380951,-0.00477328649540332
"951",0.00308581233643279,0.000256114651803419,-0.00881501650554872,-0.00411216684714311,-0.00988122699418514,-0.00289728036358372,0.00866490460075453,0.00324199551534443,-0.00249441391987992,0.00479618003680238
"952",0.00777719013036982,0.0174000528101215,0.00296428682372407,0.0184741766713226,-0.00155066530641701,0,0.00987015292083804,0.00870016627028947,0.0159896929984249,0.00477332743478698
"953",-0.00390094102814265,0.00603618132716122,0.00689658386443393,-0.00170726738376792,-0.0149441411168474,-0.00571239164989046,-0.00307664260022833,0.00689979015786113,0.00507192484893348,-0.00158359108553852
"954",0.00204331694662363,-0.00249956201956614,-0.00782755382776434,-0.00128248243584128,-0.0122157410468728,-0.00433277058813564,-0.000545225083446454,-0.00587387951178875,-0.0079406827458256,-0.0111022708620921
"955",0.00492760500090839,0.00375942481125247,0.00690335440021106,0.000428043103041675,0.00807867320772315,0.00475720679745795,-0.00508593906966315,0.00787792755313577,0.00448837545944514,0.0100240858846563
"956",-0.0131041185449501,-0.026966353394033,-0.00881501650554872,-0.0316647189990262,0.00603454722907393,0.00342493705690883,0.00492964371091453,-0.0315095295327944,-0.0310544982950141,-0.0293767432883081
"957",0.00976587202458901,0.0197586009367985,0.00790510357033058,0.015908188340785,0.00216325817900009,-0.000601835612681123,0.01998559378251,0.0214377490308288,0.0092998692698496,0.0237218936144195
"958",0.00220563877726954,-0.000503088829561738,-0.0127451684403944,0,-0.0118728465372662,-0.0055255833038701,-0.0019597092246123,-0.00864190508365037,-0.0140877695810663,-0.0123852560833844
"959",0.00186267165877219,0.000755029904796034,0.00794435517341241,0.00108753099590508,0.00675235030286814,0.000303011929722929,0.000178892976139489,0.00498111715115601,0.00200814859034404,0.0084953217711945
"960",0.00295732281149985,0.00327051565789116,0.000985300699508862,0.0108625861560256,0.00286093877204729,-0.000302920141306395,0.00196261154191957,0.00272625715787966,0.00863339269662822,0.00521452919396115
"961",0.000168316657666923,-0.00802404526185863,-0.00984264326851625,-0.000859687718766988,-0.0154422252006347,-0.00666786191593305,-0.00587676606217757,0,0.000229262503816718,0.00518756107376728
"962",-0.00286402933462038,-0.00910018007951063,-0.00298196701997733,-0.0169931369459615,-0.00879109114897514,-0.00579626910045461,-0.0100328294209073,-0.00543717018439671,-0.0103912052876222,-0.00317590168457615
"963",0.000169163783436233,0.0104593301905163,0.00299088574262241,0.00634586878823162,0.00272149288114232,0.00583006170698042,-0.00615267146159271,0.00447292565411672,0.0132798096578193,0.0051772725314605
"964",0.000760071488830949,0.000252454302498872,-0.00397608258247262,0.00282693878466667,0.00934697724069311,0.00447508875352831,0.000728689427707652,-0.000742362986287715,0.010515010266877,-0.00237718728795866
"965",0.000337714484931917,-0.00630993327788598,-0.00997990197318865,0.0110580186191671,-0.00430496751823717,-0.00167477879489042,0.00727760867465421,0.0039614588380561,-0.00527821615435886,0.0063542032704953
"966",0.00793037019369014,0.018287888519664,0.00705624647090675,0.012438184532636,0.013142890057628,0.00335497914232907,0.0056000054840708,0.0133169737508627,0.00432085361311185,0.0090765567807225
"967",0.0040176541716308,0.00698442056949089,0.00300306756332946,0.00614281876954292,-0.0203996521012171,0.0032420405024427,-0.00107780088965925,0.00219034841436572,-0.00694390493833852,0.00469301607448758
"968",0.0192582166147244,0.0240276212976667,0.0229541733145249,0.0227368918929742,0.00778392413458939,0.00807905021706512,0.0258946102106534,0.018212556831017,0.0338982424771019,0.0237446438397573
"969",0.00376246454625306,-0.0128204398815605,0.00878064664441203,-0.00185253373276706,-0.0171533387620989,-0.00420760941512333,0.0099914318460057,-0.00310037571347699,0.00257300597348387,0.00418253064980045
"970",-0.00187418073455958,-0.00833121800483783,0,-0.00412484485747955,0.00449029075213447,0.000301606513683828,-0.00485964392978122,-0.0095694503824415,0.0102653904434158,0.00265047491442716
"971",-0.00718427294794588,-0.0103779268416105,-0.00676985576205058,-0.0126320237534272,-0.022048042728066,-0.00844784953676292,-0.0361001777412538,-0.0164250388800382,-0.0158949268100952,-0.00679756808052623
"972",0.00402939505037736,0.00124807000429827,0.0116844227464841,0.00734072267861974,0.00135087002744516,0.00375283128870829,0.0119411644353851,0.00171940446351626,0.01216910575025,0.0106463598290467
"973",-0.00376769460569992,-0.00997491342132784,-0.00577473690598296,-0.00978554219560557,-0.000519339740650548,-0.00111124550070929,-0.00804585133273705,-0.0132387008504484,0.00306032486664498,-0.00827682583247247
"974",-0.011838074981842,-0.00554163971717725,-0.00774451312168412,-0.024179912392586,-0.00539775002579845,-0.00829616108433728,-0.009372565686662,-0.0134163154370347,-0.0288391826575858,-0.0417299075536764
"975",-0.0014144281631181,-0.00202601419008752,0,-0.000431114479875427,-0.0208745511820401,-0.0128529393537511,-0.0109170850612795,0,-0.00949961837834368,0.00158342810595902
"976",-0.0155792415690615,-0.0253810338169357,-0.017561035314405,-0.0262989750305163,0.0248378500748605,0.00744087326992005,-0.0314566354372043,-0.0198942585765239,-0.0109499850619239,-0.0296441914335533
"977",0.000507753828613566,0.00364590393044728,0.0148957279495485,0.0050923524302886,-0.00551284093484694,-0.00287235382870565,0.00873669717637937,0.00179892473229604,-0.00450481786283241,-0.00773932753243955
"978",0.0147181217896108,0.0238714906660824,0.0254402542654149,0.0237882970027834,0.00407879538284406,-0.00236550520825496,0.00696639932040277,0.0159011851807787,0.0131154389816137,0.0270935643193935
"979",0.00275123686171708,0.00380120901102421,0.000954471277131885,0.00064557871554638,0.00614552799889867,0.00206111712417845,0.00467462856154821,-0.00530143617106682,0.00083277313446195,-0.0143884167031987
"980",-0.000831494860865756,-0.0143903338240049,-0.00285995518268278,-0.00301012167708525,0.00424500084556279,0.00535126769814132,0.00204747555295315,-0.00380741773493931,0.00968229220156491,0.00324407562208728
"981",-0.0144768819605086,-0.033042879034166,-0.0191203323054495,-0.0317016239404607,0.0049485638707083,0.00204697399648079,-0.00705819494592597,-0.0236943009943082,0.00696739607334118,-0.00242518921933998
"982",0.0147739643033484,0.0105960062350938,0.017543715464948,0.0231624179323835,-0.0178505102077303,-0.0107250202981061,0.0192669599974034,0.0120043102265932,-0.00171126399192723,0.0186385273102563
"983",-0.0116472277087077,-0.0152030957044201,-0.0162834496697529,-0.0248148341107448,0.0138926737719289,0.00433701666677089,-0.00293624312717244,-0.0128934872421508,-0.00797430359084894,0.00477332743478698
"984",0.00303036792856792,-0.0167690713493569,0.00486868112570282,0.00781273574283659,0.00854992590798043,0.00215923777441329,-0.000552645104931915,0.00261259065774699,0.00300498833292018,0.00197938699468603
"985",-0.00562285294988873,-0.0151596875359041,-0.00484509191812876,-0.00819520655106054,0.00520983371836348,0.0017434843291948,-0.0038670003274649,-0.0122459513528781,0.0143060674970439,-0.00948249177806404
"986",0.0212679822835193,0.0321606087292703,0.0204476539823464,0.0285843893075191,-0.0222290588173375,-0.0131507072670355,0.00758005394637995,0.0269059448148827,-0.000295325657883816,0.0295174429557872
"987",0.0128085631069326,0.0229028576097698,0.00954185322628165,0.0197567589999157,-0.002607044379622,-0.00249646327644615,0.013577820568442,0.0215771368625044,-0.00132964982531958,0.00852383101731813
"988",0.00269287146336694,0.0119758810321295,0.00567114448816519,0.0036192765190064,-0.00784220102228061,0.000104546128549154,0.00144828054935076,0.0057830751477761,0.0212278850864176,0.0126777038589156
"989",-0.00105815203464343,-0.0100334359625133,0.00469945978675779,-0.00169699616921548,0.0141218415344331,0.00625669269838758,0.000542048122363026,-0.00400003906707302,0.00753236725772033,-0.00113815050425914
"990",0.000570396087831382,0.00571758008979129,-0.0121610749462612,-0.0046747704742246,-0.0214071727126377,-0.0165809530898249,0.00325207077414191,0.000251086178580939,-0.018762137741628,-0.0068363323991949
"991",0.00366337218106416,0.00594287873714539,0.00284088672235461,-0.00640498560346903,-0.00966322017958909,-0.00853516065507465,-0.0149466754887438,0.00250957207103242,-0.0125275238095237,0.00764819747851098
"992",0.00389371538458527,0.00154152740898406,0.00188869801631086,-0.00343788047202154,0.00493229763915104,0.00212620860693891,-0.0107859463823101,-0.00150193007881827,0.00430300489740354,-0.00265651027620528
"993",0.00581774703749072,0.00461588769777399,-0.0028277201867366,0.00452799812439042,-0.00608216756492186,-0.00848523433994819,0.0103492751885539,0.00350948216758384,0.000295552939925781,-0.00152208837496137
"994",0.000642701388771316,0.0104677543608735,0.0132328833740327,0.00643906379462589,0.00375768371748153,0.0032096911530195,0.00256057775345564,0.00949301151251714,0.00472637900520279,0.00990851900668721
"995",0.000883037717212876,0.00151584011902806,0.00373136772499305,0.00149281124762668,-0.0145453872778732,-0.0105563195401364,-0.010217076708083,0.00445436972989866,0.000955457531301773,-0.0026414734242225
"996",-0.00457206908826879,-0.0151361999087362,-0.00650568692627473,-0.0161842925879901,-0.0130235197755973,-0.00409449637522175,-0.0110600714780329,-0.0101012934783125,-0.010867940050489,-0.00264846928545504
"997",0.00580181788522083,0.00512294184141115,0.00561289684419397,0.00281411661671105,0.00692727471721422,0.00595158033316068,0.00260966569307719,0,-0.00660726815012469,-0.00341429533432092
"998",0.00107082482437892,-0.00713550901290183,-0.00279078403917077,0.00151136020797682,0.0182375206291394,0.00860381844228719,0.00780826912791932,-0.00971599636716725,0.00291457294543851,0.00761322130876096
"999",0.00241344529548093,0.00268695163027455,0.000932883041905974,-0.00452636270752194,-0.0010729295305949,-0.000106302308953587,0.011436986848717,0.00510755541755969,0.00678095395188438,0.00906686105773313
"1000",0.00634044738267425,0.00541074610464221,0.00591148740556346,0.014597207403608,0.00697959477128052,0.00213360195100987,0.0109427846694659,0.00909300137775526,0.00155433349452783,0.00636464767940859
"1001",0.00311055858374187,0.0035879557998304,0.00373143347736682,0.0034407598980104,-0.00714373658941636,-0.00276759531548387,0.00696587655730152,0.00715627247160588,-0.00199529992634417,0.00520837720647793
"1002",-0.00143121142750391,0,-0.000929519228247466,-0.00107162579123743,-0.00204105585881975,-0.00352184946419987,-0.00307870640509356,0.00131551118326745,-0.00288781185736087,0.00370098782268258
"1003",0.000398046844326538,-0.00689480330301528,0.00279063636530941,-0.00321809033082909,0.008931956765869,0.00385558226617522,0.00799301250461593,0.00630784523077144,0.0026733995938395,-0.0018437084596814
"1004",0.00143276014192284,-0.00128575959122235,0.00742103281126716,0.000860996329860253,-0.0195847443822403,-0.0105044670727144,0.00396481543297367,-0.000522415844552149,0.0162938596861544,0.0107130102608699
"1005",0.000714906119457348,0.00926874464673788,0.00920839508559945,0.0128026637897074,0.0169193211325562,0.0112428334271684,0.00448727004316529,0.00966813983650816,0.00357095173028021,0.00036549207135006
"1006",-0.00158811249152502,-0.00459174425523101,-0.0082117105095284,0.00509882990558874,-0.000750860991854618,-0.00203051833387324,0.00125084843973911,0.000776631768113711,-0.00493797084768133,-0.0120569444895691
"1007",0.000238681323957657,0.00666334162484317,0.0036799416883293,0.00697506704705808,0.0110642892544708,0.00503446310997591,-0.00124928577257966,0.00672314287965148,0.0123330804373718,0.0188608017722003
"1008",0.0103380316709112,0.00814676685858018,0.00916578908874444,0.00965589875491912,-0.0075439822152843,-0.00309134376972708,0.0155470164292966,0.00899040514377902,-0.00519031859003516,0.00435584443840731
"1009",-0.000551245994787619,-0.00202021658180784,0.000908307051196378,0.00457365515234143,0.00117787498535127,0.00235248388391374,-0.0177722289214076,-0.0050914499125877,-0.0235507246376812,-0.0133719597444494
"1010",0.00519779451178626,-0.00632614558361877,-0.00725951799056601,-0.00248321133699148,-0.0220273814438582,-0.0107729164471662,0.00412010174103661,-0.00230295078955145,-0.00282007421150288,0.0106226410499182
"1011",-0.00195839688641097,-0.0114590159589357,0,-0.0105808702783664,0.00437301708692206,0.0051757662841303,-0.00535224064468753,-0.0143625524877665,-0.00401870224077916,-0.013410585848192
"1012",-0.00196266894400321,-0.00540925050268526,0.00365599524298643,-0.00922623191948901,0.00533506095308667,0.00665066010002446,-0.000358775497530495,-0.00312286316171351,-0.00186804151732733,-0.00367371914114689
"1013",-0.0012586253163156,-0.00492151651300154,0,-0.0103705985319524,0.00541366657874143,0.00340981124927642,-0.000358698558319825,-0.00313238946801975,0.00404246887194981,0.0117994381284996
"1014",0.00354379509177494,0.00702760380075906,0.00728636515301262,0.0106926298005248,-0.00560026632547372,-0.00392909894820104,-0.00179526813065456,0.00418980013778869,0.00589031486319391,0.0112973335278741
"1015",0.00902491121309335,0.029465173591595,0.00904137342674782,0.0201020012017923,-0.00779801991321849,-0.00287883992848037,0.00449582998877784,0.0151237539962854,0.00407681405153615,0.0064864718915163
"1016",-0.00163355898484885,0.0047704710773524,-0.0008962032906491,-0.00871215738785525,0.00895072157631782,0.00673622597850865,0.00286426942095019,0.00154135655785259,-0.0104090058108441,-0.00143220592840976
"1017",0.00724489323427835,0.00924508241179534,0,0.0029297457076074,-0.00638366710863458,-0.00276144406144685,0.0067829839082072,0.00641201506773115,-0.0101454753417649,0.004661289919627
"1018",0.00170138814527143,0.00990354776217783,0.00269073369456829,-0.00146054273803808,-0.00468164456255238,-0.00244965753050752,0.00939742095021301,0,0.00557684067259268,-0.00107079602915094
"1019",-0.00980535615977207,-0.00833554303684969,-0.00178891301459738,-0.00773106298129878,0.00722026301244028,0.00256270915949197,-0.0119445467232635,-0.00535179367816507,0.00217348433796283,-0.00107179677897651
"1020",-0.00132572292524447,-0.00642774478293451,-0.00896035947073492,-0.0109496265808964,-0.0137933182534874,-0.00777474867145223,-0.00213311072541833,-0.0102485000774871,-0.0188453782617007,-0.0100142801895847
"1021",0.00226418963479458,0.012689683175628,-0.00994567962601434,-0.0104319554924305,0.00792920153596977,0.00332761629987832,0.0039194031903047,-0.00025901494103675,-0.00129571649304228,0.0101155804464559
"1022",0.00568687284814318,0.0100740024948678,0.00639253421929853,0.00774535456170211,0.000437232732796167,0.000106647308505403,0.00496868761723479,0.00699127115304843,-0.00511331759988787,-0.00858361088916537
"1023",0.000542276284350551,-0.00267592492361146,0.00907458946539363,-0.00597791322000607,0.00950156405419689,0.00502750876135694,0.0105949480151726,0.00539953815350613,-0.00199443846276126,-0.0126262752838782
"1024",0.00387082297677943,0.00536585323205774,-0.00179895850185285,0.0088056324075847,-0.0151464649467715,-0.00606608617733717,0.00279605474014488,0.00332504470318318,0.00814756303700692,0.0222871715082313
"1025",0.00246777101400597,0.00558003039015009,0.000900942560317697,-0.00340618888937505,0.00450408948773262,0.00374757818972671,0.0139396700707541,-0.0025488231842582,-0.0246264402370709,-0.00857762194444589
"1026",-0.0174630035188292,-0.0243669195823848,-0.0171013183456908,-0.0316174441841269,0.00524921794774524,0.00458690005896711,-0.0156381068705389,-0.0171222892638666,0.0183694129602125,0.0126171730460689
"1027",0.00751642242475747,0.014095015619636,0.000915285138898048,0.0105891816934094,-0.00761520815001282,-0.00392837339190244,0.0118710825957802,0.00832013015739386,-0.00314709858111084,0.0156639803234693
"1028",0.016008645593415,0.0246282936302997,0.0201280579830401,0.0242304991669025,-0.00495048718379909,-0.00464944551292057,0.0046584432172514,0.0180506941413208,0.00716106903677027,0.00736068056253858
"1029",-0.00191188704354361,-0.00333163669428993,0.00986569204883381,-0.00745960041254534,0.000220925559762719,-0.00236211828050115,0.000171600021685592,-0.003039559072891,-0.00267588678877939,0.00974249329415966
"1030",0.00222237209574438,-0.0050147468592926,0.00799282293625203,-0.00128836737784899,-0.00828973466551741,-0.00570486837792339,0.00257562552153345,0.0015241009859841,0.0134151018799946,-0.00654715488960811
"1031",0.00282909708476109,-0.00287945688889624,0,-0.0002150005263446,-0.0101426100350602,-0.0061702111301859,-0.00907697270794827,-0.00608820682801547,-0.00408466726364609,-0.0055498412586894
"1032",0.00625224256078494,0.00601655933351131,-0.000880995089699965,0.00129049062695463,0.00517965031668455,-0.000436386478817274,0.0112341715839273,0.0028075383156243,0.000151822872495266,-0.00279037104622348
"1033",0.00454691671057983,0.00717692088540955,0.00617286666814376,0.000429644100281568,-0.0091856361852648,-0.00686403207223418,0.00256347024531034,0.000763700163978642,0.0110875309660747,0.00664576963206298
"1034",-0.00226317250195274,0.00190053588880801,-0.00701138398845469,-0.0229716055497586,0.00870497126949954,0.00570574354156705,0.00238684222747154,-0.0094097953612462,-0.000525702272237361,0.00486435090443704
"1035",0.000378250045492301,-0.0101944759998042,-0.00088244713668284,-0.00944813956811985,-0.0115439910004453,-0.00327338552929035,0.00323123143702775,-0.00744572544016742,-0.00165327262664072,-0.00587820501003333
"1036",0.00597030958100486,-0.000478989826577791,0.000883226537411685,0.012200457562525,0.0144000783754925,0.00459763169760596,0.00627228349918796,0.000258983426713044,-0.00398945409155649,-0.00347824910264893
"1037",0.00240379436883176,0.000239625591058612,0.00882619695881148,-0.0050405659908842,0.000670630445665177,0.000326365328679579,-0.00016842993845656,0.00206849318549729,0.00476110917980832,0.00488653099623337
"1038",-0.00314773480064978,-0.00167723174446377,-0.00699929374434782,0.00198244854649809,0.00446915539619597,0.00228734495891469,-0.00336986643696913,-0.00567759694425463,0.00767208742396597,-0.0128516878535987
"1039",0.00631520248286832,0.0112794498924067,0.014096975533856,0.00835337178819962,-0.00322516892620317,-0.00141283761722277,0.00287417709425375,0.012457931007277,0.000970403814507748,0.00738913410732644
"1040",0.00298868355820447,0.00427132573032285,0.00868809210847066,0.00348808462010286,0.00156121662416231,0.00369990164328415,0.0013483479162788,0.00845961363396475,0.00700959700180781,0.00314354882990564
"1041",0.00208548796407104,0.00472607392918278,-0.000861290744263665,0.00608310935556977,-0.00311887326216154,-0.000216153754625359,0.00387224540585351,0.00279586935428844,0.00274001050933093,-0.0010444823480118
"1042",-0.0200697543017678,-0.0275166335554637,-0.0275863203571275,-0.0319585228567456,0.0149740899454953,0.00965134510101429,-0.00905598028038468,-0.0240810915513759,0.00649870005173336,-0.0013942307795789
"1043",-0.00614425718309153,-0.00096721452587023,0.00177305391106763,0.000892148731654663,0.00363327203367825,-0.00247058839833558,-0.00795393135188038,0.00545440514303119,0.0089515156112745,0.0223385505785685
"1044",-0.000686948803664489,0.00145221033438214,-0.00265473160336316,0.00245150107093295,0.00636204682767483,0.00258498073865399,-0.00545899466621524,0.000258479712790916,-0.00749035733729753,-0.00887669868527741
"1045",0.010692703498256,0.00991049671606059,0.0133097924715209,0.0120054872145008,0.00588642791180871,0.00322181343524663,0.0178389872627192,0.0178202123740492,0.00659443893887568,0.0220461048357377
"1046",0.00619655466095725,0.0117283983178151,0.00963195099306424,0.00593137173251046,0.00130059386067871,-0.00042871793921162,0.0208965520672184,0.0134486134562937,0.00203813502554451,0.00168514618857385
"1047",-0.0166728198164025,-0.0160870657256565,-0.00173450833629496,-0.010264207874334,0.00289870169280593,0.00113762103423043,-0.026906464133041,-0.0160243037884985,0.0172162932669973,0.0151413553204189
"1048",0.00213836994409733,0.00673210112158817,-0.00868806675613831,0.0136802892934682,-0.0153727827382691,-0.00525411725681779,-0.00797313487504847,0.0050890667957626,-0.00078555310137518,0.00397754323492205
"1049",0.0172242624355545,0.0128972782104735,0.0096407776599361,0.0198085992634418,-0.00978607548648502,-0.00679046473697087,0.0143641026080841,0.00860773325157527,-0.0130789167106762,-0.000330205386527171
"1050",-0.00749244443128672,-0.00848870429273918,-0.00694451023291787,0.00106722707011775,0.0083282539316254,0.00716262572335036,-0.00859767468444417,0.000501844330330847,0.00912455671300028,0.00495373116318754
"1051",-0.00785019612190463,-0.00808558575695728,-0.01923063384503,-0.0140724257617744,-0.00638731396962933,-0.00247816994431338,-0.00646148668457958,-0.00777704814619273,0.00265514879131024,-0.00460062643848858
"1052",0.00874960934580282,-0.000239549524668092,0.00445616832410511,0.013408129885776,-0.00609525098969266,-0.00237634340799764,0.0124937593129004,0.00227550031956048,-0.00257658171645725,-0.00858377702770841
"1053",-0.00143338627290623,0.000719266488265813,0,0.00192057814897373,0.00970103596290173,0.0058473360013338,0.000507191772966209,0.00327962408650739,0.000358804532442303,0.00399601803386762
"1054",-0.0185057648713418,-0.0230050748004391,-0.0248446473232273,-0.0296059375918322,0.016785915064736,0.0085043331825041,-0.0155432766383524,-0.0226302798447117,-0.0117638616522814,-0.0162520558719252
"1055",0.00692621090565626,0.00392464619390931,-0.0163785883622309,0.010316133087376,-0.00564740707507183,-0.00234771154692914,0.0113265072771489,0.00102915720688146,0.00326629155066294,-0.00573161612253437
"1056",-0.00603763168518823,-0.00464232838707812,-0.0703054853516157,0.00586576071665545,-0.000437259035774074,0.00224638449104853,-0.00678764643631113,-0.0187614200497178,0.00463029948900107,0.00271274688097622
"1057",-0.0114572684955023,-0.0252822838427609,-0.00198993855013996,-0.0166308654240269,0.0149716783825053,0.00362982653368471,-0.00803012945644865,-0.0275013353276056,-0.01865185785214,-0.0365235273160286
"1058",-0.0185128048736286,-0.0307226106711759,-0.0368892012728764,-0.0204259131448171,0.011304513897779,0.00850952513479064,-0.0130901784356816,-0.0250468003918185,-0.000220143825636065,0.00596703307699742
"1059",0.0132351140451861,0.0350740748329068,0.0455486654392516,0.012331874503454,-0.00766595418658145,-0.00305875588126403,0.00837729205064841,0.0256902591856558,0.00535816187029647,0.0310536687711132
"1060",0.00363706995580904,0.0107930143869315,0.0267328627505545,0.00177194891692345,0.00268257691488727,-0.000634977744404797,0.00882662944750567,0.0237395478242703,0.0102211724449064,0.00575298742614816
"1061",0.0154979616816413,0.0245842375708258,0.028929213418236,0.0192349585696501,-0.00588532699930988,-0.00518688535204803,0.0109794789285078,0.0237966894822226,0.00556481916473284,0.00471070698178733
"1062",-0.00346863126610508,-0.00266587494729442,-0.0037487281716182,0.0030369360936382,0.00333659319381652,0.000531743601543955,-0.00899369900748193,-0.00723131869704363,-0.000646801787025919,0.00736764965761338
"1063",0.00286182466905416,0.000728879975193886,-0.00564447062914708,0.0131919796046658,-0.00128713362088129,-0.00127601822124956,-0.00753431101168267,0.00884510428749374,0.00927718786169329,0.00199472211951734
"1064",0.00956341187956067,0.0150556322079503,0.00189234535454563,0.0115261878748609,-0.00751795146695233,-0.00511156779647715,0.0046584432172514,0.0105723659306842,-0.00798058309763683,0.0033178730098975
"1065",0.00305578546228014,-0.00885155481531097,-0.0245516000919339,-0.00105527229201852,-0.00248936763451491,-0.0026760959377734,0.00507562496380909,-0.0109719785829773,0.000287271941622924,0.00264546644963271
"1066",-0.00243707029977025,0.000724146375368218,-0.00193599994079163,-0.00506954374106328,0.00141000196163277,0.00032203090091798,0,-0.00438622787093901,-0.00517019981222888,-0.0135224126400227
"1067",0.00671859342934256,0.00410009979187298,-0.00193998173202492,0.0114648269812236,-0.00769243206471093,-0.00289779685601776,0.00448128153751282,0.00103672458543591,-0.00238188260916128,0.00568367458562014
"1068",0.00690124641709344,0.0100890587943925,0.0155489430024753,0.0128042828172299,0.00797049318180898,0.00344380968083313,0.0116675747427193,0.0111310746356692,0.00332820328993977,-0.00132973490910149
"1069",-0.00135575615338557,-0.00546966838199658,-0.0124400127009343,0.00870493753332657,-0.00205749631071805,-0.00257339301527193,0.00746283652891644,-0.000767916237635946,0.00858154624044927,0.01564586580112
"1070",0.00422351563407375,0.0119560670140131,-0.00193798893475283,0.0160262770334298,0.00486145213018596,0.00213379432362082,0.00235671564227946,0.00922345448422179,-0.00471903328529233,0.006882928416728
"1071",0.000826098655332785,0.00543474032631153,-0.0135925191764268,0.00849329819400912,0.0010843077420184,0.00225893944975386,-0.000839628519138658,-0.000253855208783182,0.00459769406460553,0.00911459275608784
"1072",-0.000149885955035955,0.00258508435159066,-0.0196848892067092,-0.00200490343215753,-0.00400966666123914,-0.00504385093118598,0.00168114577343959,0.000508129008902625,0.0158038262529698,0.00096772869811601
"1073",0.00315202664567305,0.0114864000632375,-0.00903615190274532,0.00542470286144492,-0.0150124411822802,-0.00431508406297954,-0.00134275477188828,0.00736009601031573,0.00232313969046527,0.00290047881931033
"1074",-0.00254362175724809,-0.00370777627848373,-0.00810524175292082,-0.000999192442863839,-0.00198862402946554,0.000108296195749924,-0.0104184555662296,-0.0136053474903871,0.000912979318971052,0.00192792795831886
"1075",-0.00345067066090654,0.00790860174857522,0.0194075588551847,0.00100019182697886,-0.00531245444849693,-0.00292517540595716,-0.00747132123759997,0.0107279445331034,0.00806967258682434,0.0237332348437118
"1076",-0.00301042354280068,-0.00138481625286568,-0.00701417583324315,-0.0117905001054432,0.000890311161301449,0.00130377329961617,-0.00102663488019716,-0.00732855978253588,-0.0071001320590246,-0.0184837784171399
"1077",-0.00747400023412359,-0.00970635866469993,0.00201837455214426,-0.0188071003109711,0.0107834070944948,0.00564264043618734,-0.00205494194902134,-0.00789200359362952,-0.00722096191265387,-0.020427623687187
"1078",-0.0000760277571065782,0.000933232325338595,0.00402829459595644,0.00824420842206819,0.00626828866724272,0.00388429635767129,-0.00120148924985031,0.0030789672360485,0.00204782852872087,0.00782006312591998
"1079",0.000760887545689037,0.00349729466069482,0.00702088804926482,0.0030663800652051,-0.000765781704608948,-0.00333177027710829,0.0135740335046153,0.00818629394625892,0.0134602119856329,0.00258645032519977
"1080",0.00364823274358028,-0.0023232293507981,-0.000996061848549612,0.00122272780294064,0.0135632579992597,0.00733330477286009,0.0110187661426757,0.00304521262464008,0.00862252289301879,0.00515972166490997
"1081",-0.011208656525876,-0.0251512647825558,-0.00299096127812726,-0.0250357683477999,0.00226601914133195,0.00246170141149871,-0.00989316893445924,-0.0146724822925601,0.00606680442467833,-0.00609568631687829
"1082",0.00574466981832455,0.00859982466386144,0.00299993396445197,0.0144049227939471,0.00430634830161591,0.00128120140766486,0.00779029478644855,0.0077021867964806,0,0.000322850943261122
"1083",0.0136317211742309,0.0272383186061742,0.0149551555097083,0.0236675808591733,-0.00643177674690232,-0.00394598702635096,0.0115948144340317,0.0168149891577272,0.0039060304758598,0.0158115350310737
"1084",0.00510904684810565,0.0069175126586174,0.0039296836242364,0.00884597997878767,-0.000863509269186324,0.000750728942849221,0.00714300749754782,0.0107743657900208,0.00163825938566542,0.00730619171549063
"1085",-0.00104664249255115,0.0016030755605505,-0.000978832385618356,-0.00817039189233004,0.00377962347109806,0.00353022358377975,0.00494755226731458,0,0.000885852498096806,-0.00283811777633758
"1086",0.00860519716361785,0.00983036769111223,0.000979791437208277,0.00863943427085889,0.00968249483950756,0.00426435953776449,0.0093552469950049,0.00793254677111821,-0.00333621581453702,-0.000316316289468599
"1087",0.00652869361719866,0.0178857076285446,0.0019565226763929,-0.00179272165418187,-0.0102286526579308,-0.00286611564053518,0.00455276237044666,0.0108217511390414,0.0192648715922641,0.0060107715714699
"1088",0.00324292790117986,0.00400347683178137,0.0263670646361689,-0.00818187845350715,0.00764351400734209,0.00383292321018369,0.0111686225317256,0.00389289038100293,0.00415556308623799,-0.00723270247891861
"1089",0.00235128465013701,0.00443053069223809,0.00190292653597979,0.0060361421704882,0.0030977873597986,0.00201545854707597,-0.00480216925153087,0.00484711482661515,0.0170203436180589,0.0104529163490235
"1090",-0.00153919425748661,-0.00220561096302108,0.00284905156179205,0.000199895778746129,0.00160460034784804,-0.000307938429434551,-0.0001608218614082,0.00144720263305254,-0.0128633659140043,-0.010031372377705
"1091",-0.00359716143704036,-0.0077364824315852,0,-0.0221955449386791,0.00566019471101398,0.00265377929055632,-0.00675677019130927,-0.00939273260417717,-0.00352369513932049,-0.0104496070956075
"1092",-0.00663096688148723,-0.00757410407605674,-0.00189383351944672,-0.0165642761133489,0.00445985161086693,0.00254128303591283,-0.00550690011155541,-0.0111845142542076,-0.0143448687501713,-0.0160000118565692
"1093",-0.00904801975928848,-0.0255892155553862,-0.00759009531791399,-0.00956546551995663,0.00951427853235587,0.00496325161995026,-0.00146601077095199,-0.0118023932473813,-0.0288363576480433,-0.0669918253132131
"1094",0.00441571956360143,-0.00483742084634686,0.00573642992177548,0.0130167341164678,-0.00439840412445647,0.00052580399882185,-0.00538209847550819,0.00870888525660507,0.0127552937007369,-0.00313697441194594
"1095",0.00387469541009566,0.00555528870140876,0.00380184525772487,0.00186535098711382,-0.0010515802400245,0.00147041911702472,0.00393555716751237,0.00419340008294422,0.0143152233795893,0.036713179193959
"1096",0.00853614016058701,0.0112803973302273,0.00473479104675878,0.011791523117179,-0.00716062979303489,-0.00482421883089679,0.0138843268319546,0.00245668074174632,0.00352821944876425,0.00910628911108069
"1097",-0.0105247097708262,-0.0168454399522457,-0.0169648673998856,-0.0220812792381081,0.00572783156081869,0.003582370075772,-0.0111165079408239,-0.0161726964957647,-0.00919540943321462,-0.0320855705109503
"1098",0.00476057795151119,0.00324175378630853,0.00287625484682197,0.0029271929485768,-0.00632748882212641,-0.0022052233844313,-0.000162729722941402,0.00547889504965404,0.000341224255415495,0.00103589746505772
"1099",-0.00769917528680542,-0.0159244217617729,-0.0210325534803032,-0.0218888531336439,0.00902031505785539,0.00389486232014002,-0.00912506535653668,-0.0118895785705984,-0.00654881660546602,0.00172481566061466
"1100",-0.00634135066867447,-0.000468898734655276,-0.00585936036208934,-0.0014918784469975,0.00557447239185271,0.00241057657204213,0.00230225722550492,-0.00200538579757248,-0.00178541503174445,-0.0130854680616797
"1101",-0.000150100949133036,0.00187700436495319,0.000982363576913503,0.00320165514927884,0.0102502326989746,0.00292834199904579,-0.0014766712169102,0.00728429474892445,-0.00433370036230651,0.00244246696417449
"1102",0.00893561315108959,0.00702568037328333,0.00785090952201761,0.0161701012267934,-0.0132523152126662,-0.00573494485720183,0.0111730757308213,0.00798014609128805,0.00594169524866328,0.02018793134022
"1103",0.00238183721221441,0.0083722321173938,-0.0146055522340325,-0.0064908064484257,-0.000419128880566055,0.00104826955007842,0.00194991892401064,0.0056905308202817,0.000343324161676151,-0.00784711418311368
"1104",-0.00794450096656008,-0.0161441740254583,-0.010869689331172,-0.00800822132994394,0.000524940169958077,0.00240915095703076,-0.0102171690131714,-0.00787225088189947,0.0126331004174296,0.00928471077985238
"1105",-0.0116012749683858,-0.0241444975192069,-0.0149852674749994,-0.0208200751253061,0.00482532988038908,0.00135919360966619,-0.0104866259718317,-0.017604998528169,0.00230522061478,-0.0160136901516122
"1106",-0.00083291714958833,0.00312303094444055,0.0121705935801273,0.00998043839267249,0.00375897191762742,0.00104409901872971,0.00298044671414677,0.00555296999740262,0.00514099972751136,0.0135042207483271
"1107",0.00333450092729648,0.00933897021732677,0.00200401264505401,0.00214831499198409,-0.00468109881733914,0.000103766943437833,0.00412752633410962,0.00301222203538121,-0.0000672589021404324,0.0181072403749749
"1108",0.00460763129869934,0.00972716257825046,0.0090000353376265,0.0128618390058521,0.00856988840145934,0.00552641381359531,0.0129891992080056,0.00725731802098784,-0.00242294383600838,0.00369129388523048
"1109",0.00383449382743062,0.00798885154944307,0,0.0105819733936414,-0.000414617138018158,-0.000103942824175474,0.00178541967600232,0.0111799267654531,0.00998513014448021,0.00568367458562014
"1110",0.0104111972984271,0.0219114199781567,0.0178394854948605,0.0163349521787217,0.00228058045479318,0.00155506042284559,0.0174984796049786,0.0122852603942194,-0.000400788251184836,0.00565158721344039
"1111",-0.0224608995693746,-0.0278284061173125,-0.0126582418749552,-0.0179271996072796,0.0135147681084149,0.00824096894881521,-0.0281847670905049,-0.0177186434689909,0.00180436381852678,-0.0125619145801649
"1112",-0.00106159116823679,0.00821219391523131,0.000986152341083013,0.00944205977797896,-0.019050025302089,-0.00597099017931213,-0.0057348837621799,0.00716558060168815,-0.00273500092762313,0.00870430105841091
"1113",-0.00994466154099471,0.00744683148561887,-0.00886702971466635,-0.00498870934365059,0.00574281583862901,0.00393606972120919,0.00362573085450402,0.00147213655426914,0.00481606020066883,0.00398275562528294
"1114",-0.0105812156766618,-0.015708055316261,-0.00994046793916414,-0.0160851154261329,-0.0075778682511205,-0.000619602216263893,-0.0142860042072616,-0.0100439674336067,0.00173076153820562,-0.0115702605873167
"1115",-0.000619581968460237,0.00938735065490004,0.00803223593906055,0.0078555252777881,0.00460193249390262,0.00185816009300743,0.0119939700376632,0.00296937014365106,-0.00039871080273024,0.00936459327804839
"1116",-0.00418758076569614,-0.016972759403022,-0.000996061848549612,-0.00716241663022044,0.00780996370290277,0.00216362771095469,-0.00477345698998977,-0.00764848430750731,-0.00405531184756425,0.00828362085452339
"1117",0.007631057298634,0.0130086870697388,0.00697921027927584,0.00785081068550864,-0.00402952713248972,-0.00400966602438824,-0.00926243350115519,0.00372896332364214,0.00500634143256584,0.00558665132076031
"1118",-0.0139103278869012,-0.0263832484654424,-0.00990106990852169,-0.021684194443449,0.00767577537059538,0.00320060134586186,-0.0237061426341066,-0.0173391840402503,-0.00876722248628092,-0.010457541356911
"1119",0.000783468880573235,0.00263780924009738,0,-0.00172172084223376,-0.00504422753824874,-0.0021615676473139,0.00188107710764274,0.00252079831140528,-0.00984991256198364,-0.00660506552415063
"1120",0.012686363746776,0.014111396856979,0.0199999293831081,0.0150894410181139,-0.0151062453511377,-0.00793916700569142,0.015702131869219,0.0145838590230649,0.0060905053504634,0.00698149320234909
"1121",-0.0177854635025263,-0.0360847837001776,-0.0196077752624982,-0.021447980948749,0.0181744263699679,0.0108092637438912,-0.0164676634516486,-0.0195788372518215,0.00302681782507319,-0.0267415394978376
"1122",0.00220439458625932,-0.000489595542497612,-0.00299984642285034,-0.00759568679603473,0.00453986170273235,0.00277618124722379,0.00700480332213904,0.000505569836483311,-0.00100586108522871,-0.00407053551353975
"1123",0.00298421488308698,0.0124849193302385,0.00300887257849181,0.0013120328047449,-0.00472444079434609,-0.000717530022156687,0.00848301059913537,0.00319184270358042,0.00651138479887625,-0.00442780233597684
"1124",0.00511621396812112,-0.00362682709973527,0.00100004607606285,-0.00152869479126261,0.00123833252634453,-0.00153925811326072,0.010599293573222,-0.00254516922252035,0.000600220080029246,-0.00547389412708488
"1125",0.0137037612819033,0.0232683309081294,0.0169829241703781,0.018372743785275,-0.00443220822885082,-0.00133626593631819,0.00882276407744009,0.0130135503897404,0.00486566689905787,0.000688055927610343
"1126",-0.00602544605854738,-0.0126057234036142,-0.00118894915360535,-0.0099569181091631,0.000620995789684553,-0.000411365865016555,-0.00214506005232795,-0.00881617528579737,0.00152566998957515,0.00446882846379237
"1127",-0.00287556480315643,-0.0122760075884117,-0.00198425641296007,-0.00131452952297328,0.00765683147733598,0.00525091084030915,-0.0183563452596158,-0.00304963630487953,-0.0175508902062754,-0.021218265704642
"1128",-0.0116134961916081,-0.0156601792052573,0.00596420196315517,-0.00175535783294978,-0.00421014084078775,0.00419902260967042,-0.00108776691327128,-0.00994115338671475,-0.0140218488343495,-0.0118882007975992
"1129",0.00891109996757788,0.0111112142332213,-0.00494067714318525,0.0116484031272548,-0.0137140299574968,-0.00387559666941861,0.00527561178349334,0.00437688408350412,-0.00362367713741552,-0.000353779382827213
"1130",0.0130529936466399,0.0119879362640076,0.0119164432720176,0.0136866788061656,-0.00805027696998972,-0.00921484169528874,0.00829534525429132,0.0125606529436333,0.00349968444382576,0.0176990911858448
"1131",0.00856417511566465,0.019496713679064,0.0157019015425761,0.00921554123988466,-0.00663984002794038,-0.005993536085383,0.0110812023106164,0.0091140041476836,0.00642770765769596,0.0180869597716493
"1132",0.00956230317956086,0.018639503926573,0.00772938599115847,0.0108304867238247,-0.00159121584609312,-0.00343119483928722,0.00132839848475985,0.013045589129884,-0.00801734648811947,-0.0105910798016576
"1133",0.0147758713918189,0.00879267925761185,0.00862908877616864,0.0117646900469017,-0.00159981128043418,-0.00249845100670087,0.0179105690231245,0.00841996180313953,-0.00732881506849314,0.0013812676985363
"1134",-0.000820784852727852,-0.00777377040453753,0.00190118214107526,-0.000415273771317226,0.00224237849756204,0.00628951828681812,0.00619087327152323,-0.00736760386393709,0.0186297669937789,0.0134482335920072
"1135",0.0011953386775676,-0.0104463777163839,0.00569236671850049,-0.00664726628226664,0.00511588423346554,0.00177129738973569,0.0061526226153108,-0.00395817079656979,0.00867031739245672,-0.000340247139329009
"1136",0.0103756076859811,0.00791738334906356,0.00660408258928058,0.0138018489831744,-0.00296900255224886,-0.00384747133369079,0.0125527660167548,0.00596153115956533,0.00161164457426244,0.0211027479228436
"1137",-0.00709248632909254,-0.0147583028205247,-0.00843529105848029,-0.0113451214835576,0.0141426450261182,0.0106476308838535,-0.00349673748736212,-0.0069137894314838,0.00737516623701651,-0.000999986380040063
"1138",-0.0180802231904671,-0.0374486206165149,-0.0122871142259852,-0.0279572394566919,0.0149945119566834,0.00764432584922869,-0.0188199056943552,-0.0236200602803999,0.00891844259567387,-0.00767430506191968
"1139",-0.00431916317873626,-0.00803220784761505,0.00287062711595176,-0.0100881547873406,0.00340912724987907,0.00143515263181082,0.00341377246812113,-0.00127339704356388,0.0077842076069452,0.00874238413852768
"1140",0.00334843006347207,0.0156881318877908,0.0190840596505772,0.0162619560620985,0.00277943015551219,0.00163752611909684,-0.00842394557860371,0.0104540098928709,0.00896769630247563,0.0136667549848453
"1141",-0.00690217440979013,-0.00722486925089005,-0.00936342055880346,-0.0106676867930389,-0.0142705879855071,-0.00572312163265198,-0.0111093148643284,-0.00782215459406888,0.00259500455816153,-0.00559029126745914
"1142",0.00580477206211127,0.00150585305172402,0.0075618500140251,0.00625388722053022,0.00166623695734236,0.00411180498155073,0.0109037193962738,0.00508641287546885,0.0042707650439715,0.00892861944212275
"1143",-0.00820120307299321,-0.0175393753697389,-0.0121955223907328,-0.0115730757721589,-0.00967039929403368,-0.000613912297860009,-0.00898808045757282,-0.0129048834607496,0.00882738419125095,-0.00557203579296839
"1144",0.0162315728280591,0.0132617981471002,0.0123460894004541,0.0145274651922966,0.0207899679122128,0.0037896366919834,0.0173151633675781,0.0115353854721298,-0.0121990350297424,0.00692156308141456
"1145",-0.00060256893884969,0.0135918769992827,0.0103187120326502,0.00299200418421219,-0.0118288379216406,-0.00489814390890286,0.00745650701801392,0.00608218849594477,0.00879348225026555,0.00327327776015629
"1146",0.0138709901051031,0.0273155805435226,0.0083565681822797,0.0159812779071986,-0.00770318056114061,-0.00553743174589461,0.00643614034898565,0.0118387223725065,-0.00762723990187819,-0.00489389755420977
"1147",0.000669120643106202,0.000483497940911626,0.00184166099932415,-0.00062913085802685,0.00755331273008264,0.00381495225222128,0.00511572850590092,-0.000995781077172797,0.00833167334067442,0.00819671052420667
"1148",-0.0055727360156701,-0.00579844973888288,-0.00367655103798981,-0.00209864291462192,-0.0109320516619047,-0.00318466611973744,-0.0112930731553041,-0.00647882778197728,0.00781450832098751,-0.00487801563658707
"1149",-0.00373625880766837,0.0068041178744187,0.00184505897247522,0.00336488528208512,0.00684197058387359,0.00422586388526947,0,0.00476512532346729,0.00273298595990812,0.00784313079179988
"1150",-0.0204754618516355,-0.0263091885743247,-0.0165746559818115,-0.0176064865488316,0.000104476371926232,-0.00164230436839874,-0.0268660163618237,-0.0154762677235921,-0.00367625014448247,-0.00680941221417808
"1151",-0.00290972415512292,-0.00421440816425078,-0.00187237532666229,0.000853535650143789,0.00376337605369903,0.00195308349754164,-0.00148803355753291,0,0.000827056418003069,-0.00326472866915961
"1152",-0.00683456100243429,-0.00199118428134104,0.00469009915235796,0.00426339449077884,0.0197879517639077,0.0121052164330107,0.000496828059569632,0.000253287203852759,0.00616568749580604,-0.00818865621833109
"1153",-0.00425279460171002,-0.0164630741595551,-0.00933711189194986,-0.000848879400156988,0.0100921870214588,0.00363762685669622,-0.0132385427355001,-0.00481606154460923,-0.00360093515197779,0
"1154",-0.0255474593797844,-0.0304338646853882,-0.00848228744747481,-0.0308052324056129,0.0300264811695843,0.00921230505488535,-0.0293480044867909,-0.019103722698692,0.0240933488201032,0
"1155",0.00541885569306189,0.00706272107627548,0.00190118214107526,-0.0035073459260262,0.00196976339521915,0.000802349717177409,-0.00621934690861947,0.0111663096772299,-0.000185729316846794,-0.014861261469488
"1156",-0.0468416553735269,-0.0727271960636091,-0.0607210667849999,-0.0571931190643828,0.0355808278694769,0.013230282178315,-0.0483309670728588,-0.0606063053058453,-0.0052635207980829,-0.0378813261809202
"1157",-0.0014966616985489,0.0240895390918121,0.00909069790648354,-0.00653290303193721,-0.0288531951497673,-0.0115742951823562,-0.0206430232683138,-0.00328048029366645,0.00690986682588313,0.00418112739105347
"1158",-0.0651235763319351,-0.0820569112783894,-0.0480479168273795,-0.083372616480161,0.0315673730948962,0.0159133836958487,-0.0850591779100859,-0.0811850013429679,0.0331993508500772,-0.0371269529125423
"1159",0.0464995942722632,0.0694276981734936,0.0515247106707739,0.0586727514800249,0.0030318004909593,0.00581186392417177,0.092558905480322,0.0799999114309353,0.00891578533137238,0.00972978201500774
"1160",-0.0441778933534699,-0.0696571951600999,-0.0460000500459308,-0.0530009312005489,0.0297534863940492,0.0132222757135148,-0.0235119035344261,-0.0527913921130917,0.0354071583215281,0.00428252295001075
"1161",0.0448838638152782,0.0488170086582729,0.0377359777869584,0.0552009896628576,-0.0504496619165935,-0.0146926710003343,0.0466272801571515,0.0469799447211732,-0.0219383775697288,0.0216773984576242
"1162",0.00673335346525894,0.0251287297816032,-0.00909116543426836,-0.000484719961503455,0.0198031446559963,0.00696521975189168,-0.00146068632465446,0.007803713053393,-0.00456807613469989,-0.00139135691917081
"1163",0.0211644868500138,0.0239551901784598,0.0122329507544976,0.0232615551461473,-0.0101356542064377,-0.00370175552593699,0.0356555010015787,0.0210176197922187,0.0107666175750627,0.0121908874330814
"1164",-0.00853881534564915,-0.0174101901435993,-0.00805662623670911,-0.00852474052038477,0.0165554445565539,0.00459555904241471,-0.00370742440805671,-0.00839618592784985,0.0123399008322485,0
"1165",0.000669007925972132,0.00664445842761396,0.00101501553977301,0.00716479948279769,0.0175088217673487,0.00700864132310119,0.00124041516648976,0.00655549446827286,0.00287488503765965,0.00860291493408494
"1166",-0.0431186010604724,-0.0539054023269565,-0.034482635194412,-0.0471893508892496,0.0205388469310472,0.00522057127821984,-0.0430091473087292,-0.033107272244328,0.0189198660580194,-0.0245650104809031
"1167",-0.0163306273805073,-0.020058116049377,-0.00945392699923453,-0.0124444311529371,0.00806738613546854,0.00105749345388406,-0.0199740640933549,-0.0117879736989015,0.0125478054661952,0.0178383776501641
"1168",0.000799152452734209,0.011569216606202,0.00212081465124792,-0.00100795226659778,-0.00251756746848042,-0.00182518122428466,0.00188705822367652,0.00369225056505118,0.025784935133953,0.00171818966189541
"1169",0.0329105687243765,0.0340177556203636,0.0190477939730282,0.0350656234094286,-0.013794031807128,-0.00404197103867099,0.0246753070432282,0.0271650885139418,-0.0374884779779724,0.0102917024523768
"1170",0.0140843031816751,0.00425408756265466,-0.0114225869943061,-0.00974917358124638,-0.0284300075937584,-0.0107256582827442,0.0112134218949482,-0.00110243106996089,-0.033883064489031,-0.0101868622966957
"1171",-0.0152441230003013,-0.0276760213619156,-0.0136554562479468,-0.0194434788704221,0.0108206044177146,0.00615342988296974,-0.0210872110736438,-0.0170984243279065,0.00413636484018753,0.0044597718600301
"1172",0.0145342443406817,0.0116180626224636,0.0212992569867578,0.0170682803735136,0.00986699904722976,0.00320390909455037,0.0148558911113847,0.0134677805397374,0.029647249769974,0.0112705134484055
"1173",0.0287360566700758,0.0267009561591574,0.0135557511055189,0.0323295149340619,-0.0138268534817001,-0.00658031311687968,0.0318391523985007,0.0271318277625823,-0.0201724346640422,0.00337722592734591
"1174",0.00263691345139616,-0.00782975635718064,-0.00411528647304493,0.00143437641906319,0.0160772349779792,0.00691534360522406,0.00390148827608727,0,0.0299615103223965,0.0134635385750419
"1175",0.00443751663022507,0.0194474025949782,0.0175621589813106,0.0205300823389594,-0.0154542213948486,-0.00357873200645464,0.010775684293578,0.015094320432639,-0.00770522028904908,0.00166055506291896
"1176",-0.0104723837304506,-0.0102295400850394,-0.00913731315010624,-0.00538006138922131,0.0211982194436617,0.0079689748406444,-0.0167777950573361,-0.00929395232841645,0.000843990542178652,-0.00696293982860552
"1177",-0.0255503716458777,-0.0270948014783943,-0.0163933585629896,-0.0225775083409199,0.0324859106872657,0.00917078053920939,-0.0241732495666658,-0.0144730503564647,0.0301906457016543,-0.0053421641792456
"1178",-0.00729734705239493,-0.0422050546898937,-0.0218749066799118,-0.0103467642048435,0.0103987662864886,0.00133913711121947,-0.00218558468531649,-0.0190375963880636,-0.00185555004760019,-0.00335688875632811
"1179",0.0282076491334471,0.030575604053805,0.0191690386164234,0.0296621673275199,-0.0190886370624945,-0.0053502454754969,0.0335884869577761,0.0202389439546462,-0.0318206243352855,0.00909395082323083
"1180",-0.0103914237933299,-0.0206517331026982,-0.0125391295190028,-0.0221960942149679,0.00896808066215571,0.00489879355831269,-0.00724133342377131,-0.018750002190943,0.0267110681419576,-0.00667547638088173
"1181",-0.0262099464288824,-0.0380159182938418,-0.0232802935440781,-0.033808258761873,0.0106652537165781,0.00487414199905278,-0.028108560356034,-0.0288011258354386,-0.00610528030477187,-0.0157930705888282
"1182",0.00646996371046682,-0.0101882628607262,0.00975068142880531,-0.00199927739582595,0.00105541994900848,-0.0030435115339299,0.00311169351337992,-0.00228067635220341,-0.0223021531096097,-0.0023899317720053
"1183",0.00917135948268011,0.00842162767284127,0.0171674188746163,0.00150274949541007,-0.0142320591280859,-0.00295721256460424,0.000912544801320525,-0.00343024019976801,0.0105846777674159,-0.00308004014999508
"1184",0.013843769478618,0.0238168260655915,0.00421959366068902,-0.00275108315567285,0.00846674910145695,0.000574482460217185,0.0056518649149695,-0.00372792880615092,-0.0074492329570105,-0.00480608216168577
"1185",0.0172575297246809,0.0259819708321369,0.011554570076183,0.014543633355399,-0.0152885972096178,-0.00745965390740722,0.0193980726423182,0.0146803296699931,-0.0158569656847878,0.00413940847517402
"1186",0.00591838561259639,-0.0029445217050923,0.0103839324076662,0.00173003815686812,0.0072694621599525,0.00192703060141541,0.00818044262227313,0.0000858646125032614,0.00934635926650329,-0.00446586426941942
"1187",-0.00995689683082079,-0.0318962296788426,-0.0143881538254976,-0.0296073562207441,0.0190659736569152,0.00817342154174061,-0.0197565675909636,-0.0234685300508576,-0.0154519173746062,-0.0169082305750911
"1188",-0.00116396926220463,0.00671151096731126,-0.00104265494911338,-0.00737344387295469,0.00419667671880752,0.0013359955256067,-0.00287918938953702,-0.00175869320279542,0.014251924461969,-0.00175497785306811
"1189",-0.0294581487800003,-0.0300001951959137,-0.0125263075982663,-0.0371418511355177,0.0330838433728484,0.00428656751309386,-0.0478253190097503,-0.025836717303435,-0.0124587723999247,-0.014767839573728
"1190",-0.032324411105197,-0.0390501042435322,-0.0158563703862786,-0.0702311911846395,0.0375866675420924,0.00929482691655048,-0.0252083758813954,-0.0334539188494462,-0.0261535405531089,-0.0353319713791268
"1191",0.0060252670600045,0.0117033837898504,0.00322250587413642,0.0266096143500165,-0.0185995684539099,-0.00826986001826635,0.00803840724116078,0.00904280358706067,-0.054717538218559,-0.0177581084843996
"1192",0.0237800623546915,0.0285988950180329,0.00535340530983963,0.0150498513185011,-0.0160558465022607,-0.00416946099550508,0.0126730872674197,0.0117429365371935,-0.0138923714538353,0.00338990068006195
"1193",0.0111836870459694,0.0296782885722571,0.0159743580193252,0.0318508026969739,-0.0153085876860302,-0.00666124256185319,0.0105890003043478,0.018631663557289,0.0193552669202277,0.0168919313092548
"1194",-0.0204184697222836,-0.018203740615875,0,-0.0300692344769604,-0.000341347908511036,0.000191888506407611,-0.0249569462157249,-0.0194904705598089,-0.0274544223540304,-0.0269472233298083
"1195",0.00790346002948317,0.0222496495543847,0.0178196417841365,0.0137175006940651,0.00692128572418582,0,0.0148494960415051,0.0149849635709332,0.00947379330768272,0.0117601987558278
"1196",-0.0249892553343501,-0.0365780531759462,-0.0257466224064866,-0.0500679225895135,0.0251187166816362,0.00632135375295029,-0.0263767719549458,-0.0343478689436033,0.00228282185699724,-0.0344957184688444
"1197",-0.028457784042953,-0.0313774271194351,-0.0158563703862786,-0.0210824623997574,0.0275199229081076,0.00926040872165035,-0.0470634634184159,-0.019032983989714,0.0183475201612997,-0.00504847487959281
"1198",0.0219228025108014,0.0223517698157314,0.0128894641955548,0.0154250850590902,-0.0126806596401796,-0.00510273048846954,0.0377671046034824,0.0104964800603173,-0.0206262913495028,-0.001951653922452
"1199",0.0185153848309791,0.0186947334635035,-0.00424162930249594,0.0232157510814019,-0.0071988922214139,-0.00417871741825404,-0.00759821789025372,0.00629522053419351,0.0115453438946038,0.0140790482234632
"1200",0.0180912826900705,0.0339034057429874,0.00425969735963627,0.0330532090716482,-0.0184576503468351,-0.00696280983530095,0.0276041543599288,0.0272131655811345,0.00645928731208456,0.0208252518572627
"1201",-0.00669578031652207,-0.00842365994926619,-0.00530231271993964,-0.0119307630855507,-0.00738728900404606,-0.00518601429593946,-0.0282352677082112,-0.0024360138180457,-0.00816257685330624,-0.00453344997004712
"1202",0.0334456357020512,0.0445993871289514,0.0255865172211065,0.0447310028124863,-0.0141237680965781,-0.0105230841754795,0.0482243274936041,0.0335777035824913,0.0256942529203403,0.0223909381486429
"1203",0.00100350819743533,0.0002906288472726,-0.00831600994146675,0.000525527740196097,-0.00334584055849063,0.00331732352244818,-0.0184793973065864,-0.00797436851253019,-0.00716603155102513,0.00742391804903431
"1204",0.0087718165187991,0.0223576654815372,0.00628929425415103,0.028091476821499,-0.0145464480438889,-0.00340414035619985,0.0162779538159619,0.0214352227888961,0.00715600837177011,0.00184234981324116
"1205",-0.00198749041283797,-0.00198811681386857,0,-0.00893775169338573,0.00995714283601234,0.00400107737075039,-0.00694735237413746,0.00466319363363299,-0.00588014228470357,0.00220658761071491
"1206",0.0170940819887095,0.0133751385486396,0.00208334883959749,0.0200979301807567,-0.0145293187313909,-0.00495696354402375,0.0231249941133811,0.0165359942384478,0.00677751681865324,0.0227523610500662
"1207",-0.0190912826375641,-0.0292051515213624,-0.00415782454483804,-0.0338469885263394,0.0172885417842397,0.00654421068021205,-0.0229822363422271,-0.023116253255955,-0.00477355586683803,-0.0143524120639776
"1208",0.01954585024987,0.0161988942904028,0.00939447402815707,0.0266668390165714,-0.00621063280299206,-0.00106700329058507,0.0330482813025519,0.00964056112082967,-0.00479645199841494,0.00546057776377684
"1209",-0.0118289165843256,-0.0170793585284169,-0.015511901669925,-0.0190987022401998,-0.000347349325238611,0.00155405222700766,-0.0124201790187366,-0.0144676930302475,-0.0121725225450452,-0.019551117232251
"1210",0.0043757359162111,-0.000868721962485774,-0.00315154196560985,-0.0192108078458827,-0.00712057012489398,-0.00203679616371766,0.00609765402353246,-0.00411050308616201,-0.013135616849178,-0.00147700870732781
"1211",0.0189871394069761,0.0315941202585952,0.0105377016414687,0.0285865351331644,-0.0105823911400461,-0.00184672723845247,0.029545596027678,0.0250593912642778,0.0110920958080218,0.00517744365051964
"1212",0.0122609322202518,0.012643891397299,0.0104272131222312,0.0391146736449026,0.00167966349647597,-0.000486860586854099,0.0264900416221683,0.013229796660267,0.00940320939309913,0.0158204292876116
"1213",-0.0194439887074269,-0.017480470572838,-0.0144476666600988,-0.0198117972960954,0.0254142035372138,0.00857244534426216,-0.0154125416330542,-0.0218565858438923,0.0283815171188295,0.0032597558763543
"1214",0.0101587085361934,0.0180741326572116,0.00209404437180982,0.0184439489838706,-0.0174693597489309,-0.00734049401465997,0.00928328151716751,0.0078352934050494,0.0109305999379332,-0.00577620555844283
"1215",0.0348352948690669,0.0590844631659644,0.0386627669194077,0.0607786486128963,-0.033897565585547,-0.0120654281148754,0.0427412909589908,0.0457814971614527,0.0128435428737232,0.0265069102104287
"1216",-0.000233354117923246,-0.0125718454948762,0.00402420360203104,-0.00841896580731272,0.0105175132573925,0.00600776677097303,0.00311297089754969,-0.000825774369188625,0.000412810373114469,-0.0042447971617956
"1217",-0.0241058180258461,-0.049867677365294,-0.0581163671145032,-0.037500047399771,0.0396552471974208,0.0134127151475458,-0.0131034984053013,-0.0338932740612079,-0.0134418056078823,-0.0152752847674487
"1218",-0.0278883666401574,-0.0424342940696935,-0.0127659294221225,-0.0242584940690308,0.0334740886399794,0.0119941796185461,-0.0337177001952104,-0.0199660208315005,0.000239088089855066,-0.0119047844473724
"1219",0.0163113859098218,0.0134109609792838,0.00323257998218796,0.0306375303599331,-0.012473805074286,-0.00239136034935628,0.0202499475102274,0.00407438010070815,0.0100369993417075,0.00620655986768326
"1220",0.0182272364752323,0.0322209682486647,0.00751880750565781,0.0102340305263866,-0.0137334680229906,-0.00469823550710335,0.0113410839201658,0.0133331505036163,0.0157340768453103,0.0123368135976034
"1221",-0.00609876017321687,-0.0167223493155276,-0.00213211981727557,-0.00651225309926606,0.00120359187563701,0.00298649452901367,-0.00753467069414504,-0.00514898976830802,-0.00506635799518773,0.00322572541378996
"1222",0.00621598429421422,0.00113391777240901,0.00854713454957623,0.0084971483938141,0.0063527478682992,0.0011522996654072,0.0024718795271943,0.00373820918963474,0.0241731920103063,0.0146481467086375
"1223",0.012830704230768,0.018119892435855,-0.00423735007357562,0.0117959344289469,-0.0127963804950388,-0.00450899854916365,0.0119756789400303,0.0117442541484596,-0.00828664437733784,0.00492958259453546
"1224",-0.036909627561714,-0.0631256185084377,-0.018085102585241,-0.0585299543622672,0.020740156356704,0.00886665764618977,-0.0449005414557971,-0.0450164839804162,-0.0084134847485362,-0.0220743406300569
"1225",0.00941871054911769,0.0175126702497044,-0.00108332198767846,0.00657086622893277,-0.0148999952079761,-0.00487217486809388,0.000911080590052293,0.00326082372769387,-0.00540482339842074,-0.0010748689279797
"1226",0.0188222523281669,0.0306299636577279,0.0108457528590291,0.0241024516800823,-0.00610211499083213,-0.0046078367973198,0.0258510855786052,0.0260047779289776,0.0164777843664707,0.00968441420898558
"1227",-0.00947420119838849,-0.0209451446821777,-0.00429169176423405,-0.0137287481179347,0.0160829202508774,0.0062693770051605,-0.0200534775549414,-0.0207374956177951,-0.00436887772716632,-0.0106571575633633
"1228",0.00494164623052185,-0.00578219629296217,0,0.00621431866089517,-0.00136155182751352,-0.00134234730727256,0.00869287577599698,0,0.000923810639557932,0.00718126704142441
"1229",-0.0158629778248781,-0.018028500927582,-0.0183190546685358,-0.0269269417121717,0.00911811471726409,0.00364736110667363,-0.00951525363878636,-0.026764762041125,-0.0106714697123242,-0.00249550960909894
"1230",-0.0158765346099495,-0.0106604648837501,0.00109765545279017,-0.0253870854199474,0.00802248329414867,0.00200743835689043,-0.0179445442571117,-0.0163188553970252,-0.0257127230398438,-0.0232309291562415
"1231",-0.001064798249096,0.00329253580453881,0.00438602974272162,0.00390690241784508,-0.0002514204305748,-0.00372155147496156,0.00719808776935094,0.0061442682653603,0.00311184309592405,-0.00146353550983858
"1232",-0.0190193573129206,-0.0256563034999496,-0.0196511494935859,-0.0321742365023518,0.00594876747268613,0.00277788212776597,-0.0263881798962712,-0.0262592990551541,-0.0245793767026421,-0.00732866692535983
"1233",-0.00392795685781111,-0.009798015099312,0.00779546853298241,0.00348531226407944,0.0111624520887832,0.00305609064858081,-0.00282329590181041,0.00689838771668305,0.0110703241590215,0.00664450312592546
"1234",-0.0220655194957972,-0.0303028368185133,-0.0232041652647367,-0.0323268245850867,0.00980305395223269,0.003428295773787,-0.0294451107975544,-0.027717129183745,-0.00290361143189899,-0.0150348950280789
"1235",-0.0018876531939388,-0.00510221512732278,0,-0.00331328436722333,-0.0145211043777905,-0.00635806460026866,0.00350107865823346,-0.000640617384381814,-0.00867565359854827,-0.00819058292561925
"1236",0.0289671037667631,0.0503206226850306,0.0282807348530085,0.0479227503059938,-0.000496639938219912,0.0000955740531014548,0.0244179713872568,0.0326922250429482,0.0197675099057839,0.012387333873749
"1237",0.00283994033371071,0.00640816794814314,0.004400248853204,-0.0044939491527255,-0.00819942866836332,-0.00191014836532699,-0.00283769102903897,0.00682803358356998,0.0015003300275962,0.0129774726077585
"1238",0.0411496064770551,0.0527593187373685,0.0328585694003778,0.0624002784707554,-0.0156158182555906,-0.00583666281777628,0.0461013898226514,0.0554871184468333,0.0194750713244525,0.0117129078004778
"1239",-0.000159585777221083,-0.00576054754133992,-0.0137857860630138,-0.00299924845056754,-0.00501758562226928,-0.000289634307428122,-0.0101558126507894,-0.0175232907081708,-0.00293892896787962,-0.00361785859813823
"1240",-0.000880377507101793,-0.00144833984919468,0.00322587729230239,-0.00300827100271139,0.0140170229657899,0.00443705328951238,0.00164918877182862,-0.00356714763590893,0.00112009664799562,0.00871458986637008
"1241",0.0108918656955734,0.0104440537888983,0.00750265772806435,0.0163441557963899,-0.00202284351724646,-0.000576096019820449,0.00932853848803927,0.0137231530605906,-0.0147214691847233,-0.00539956831462385
"1242",0.000317142971465678,-0.000574097440857235,-0.0117022917480404,-0.0136071697068467,-0.00954349324020742,-0.00259430573594144,-0.000725128952759224,-0.00706309820213413,0.00513976789398529,0.00542888193349578
"1243",0.00372248820592969,0.00660712550904541,0.0139936324130381,0.00401301931478915,0.00358121281237334,0.00452771299382704,0.00943056164253431,0.00533474479085294,0.00725413872505043,-0.00863930189363515
"1244",-0.0219365035149706,-0.034246636267711,-0.0244162735193584,-0.0359729350314039,0.0124903656240758,0.00508365608281602,-0.0238950554015259,-0.0341977773861811,-0.0201888909157812,-0.0127087255023969
"1245",0.0169421845865148,0.025709387145767,0.0228511472853616,0.0202122866022627,-0.0205605381017966,-0.00687031134191252,0.0198787690609932,0.0149571238126442,0.00253041336378867,0.00367777219365739
"1246",-0.0145971067014713,-0.0342842050625116,-0.017021249487754,-0.037592002269499,0.0111391124051765,0.00345857422910711,-0.0178670220229072,-0.0315787292976352,-0.0265023386959977,-0.0128252236904338
"1247",-0.00933938866509065,-0.016706513079113,-0.00432906775752595,-0.00923713742603682,0.00932094399012806,0.00459620394240079,-0.00881979399068034,-0.0102485329546853,-0.021853249526105,0.00408313009436156
"1248",-0.0106459775622657,-0.0109224886605617,-0.0108693006794185,-0.0143847739038695,0.0188895878791979,0.00419294411527793,0.00574664549210135,-0.0128651104381142,-0.0350899217751327,-0.0354898435017028
"1249",0.00361444255333043,0.00429477615567242,-0.00219810416138699,0.00648648217728498,-0.00370768601369986,-0.000854184543026437,0.0136404540466513,0.00985397403147381,-0.00366274448075565,-0.00498276289883115
"1250",0.00148253740612092,-0.00763592780927846,-0.00330406924794935,0.00751883531188802,0.011661412011911,0.00484476717048388,0.00836548008799087,-0.00331912797469647,0.0190375760646284,0.00808941651852191
"1251",-0.0106916480960298,-0.0044757579665119,-0.0143644467277372,-0.0258528550473527,0.0126723537441207,0.00340367288381827,-0.00973857222547514,-0.0150495383328703,-0.00231914584343618,-0.00458549768908145
"1252",0.0302600247952658,0.0384014270795721,0.0256409034018072,0.0419025221639535,-0.0249460657195374,-0.00904499902501477,0.0302310184011025,0.0367361479680481,0.0136243369801878,0.0230327116103957
"1253",0.00193688715927309,-0.0054117022115332,-0.00995572972158199,0.00318128812392859,-0.0139091508059495,-0.00323275373154364,0.00141452501070494,-0.0119161811199424,0.00114669387556865,0.00712943567986613
"1254",0.00885853058790453,0.0120919153515384,0.00670388467158078,0.0132137536828851,0.00419803444166167,0.00124016914421765,0.0136808892778402,0.0111077160918112,-0.00712656510240339,0.00111779615846253
"1255",0.00894085270873246,0.00567487446306503,0.00776918426721851,0.00391220962500327,-0.0111207463341721,-0.00409597300133813,0.00492696202746234,0.00784668123746779,0.00173035767823948,0.00483808137586306
"1256",0.000791009792873831,-0.00267297813559586,-0.0121145166426762,-0.0096130107394149,0.00475026119186639,0.000565236322784157,0.0022763304090283,-0.00653997823345376,-0.00895652241003819,0.00444445986150788
"1257",-0.0131231860773839,-0.0157832377392624,-0.0122632053712386,-0.0167891075947301,0.0184891654630814,0.0063213524132173,-0.0108318015156272,-0.0163008389480789,-0.0250468329985969,-0.0117995140293872
"1258",0.0103339150205788,0.0160363431557582,0.020316079013817,0.0114729864280889,0.00182336186566912,0.00123734336623205,0.00830123236556557,0.0114723031879587,-0.00456864864310824,0.0029851108523391
"1259",-0.00491605798506545,0.00476478642334022,0.00774333831233132,0.000791241167787282,0.00322681652566592,0.00351666038794085,-0.0049049095546847,0.00283547106513393,0.0109751832107272,-0.00148807495388825
"1260",0.0159362756079462,0.03141670499283,0.0197583060943645,0.0305745832249238,-0.0150102271566781,-0.00634599392894908,0.00616104243915139,0.0248192462377828,0.0258569173676915,0.0298061975373973
"1261",0.00156861078151116,-0.0103448798336412,-0.00107608902975964,-0.0056265647869852,-0.0118898147477703,-0.00314594516811018,-0.0111966093681868,-0.00367836369667029,0.00506675865914263,0.0075978046715317
"1262",0.0026623864748434,-0.0185829967405837,-0.0118535501756563,-0.00437280342750768,-0.00177945978842364,0.000191448084585044,0.00725417627375702,-0.0101540706761304,0.006827847311627,-0.0136445958527361
"1263",-0.0025773162099304,-0.0121303572224879,-0.0109049482362991,-0.0126578147625653,0.00789452481505926,0.00392007163900066,-0.00175652808113413,-0.00590603738773765,-0.00367601726249223,0.00436834231689986
"1264",0.00242757125896764,0.00509147837249246,0.00330773595659561,0.010465493283855,-0.00176858528140544,0.000189891105762507,-0.00281539994325175,0.00250120242059415,-0.00445290720966107,0.00108748494039279
"1265",0.00867063052176742,0.0146009003817038,0.0120876994213459,0.021750405306987,-0.00168707174170202,-0.00199968262668004,0.011116865971438,0.0155960569717657,0.0136741150159743,0.0072410675824528
"1266",0.00054183881414116,-0.00616760749849887,-0.00434320193413862,0.000760403938078413,0.0130151842905455,0.0058202490996051,0.00890044579203719,-0.00061434354197365,0.00649268158404359,-0.00287566377870796
"1267",0.00239936328440771,0.010047391988864,-0.00436192941967273,0.00405183009584742,-0.00141844772549204,-0.00208659526550847,-0.00657287304624943,0.0129070620517204,0.00444671515559247,-0.014059040274147
"1268",-0.0051733871470182,-0.0184317735225036,0.00219030044332302,-0.00907942765770653,0.00994186599584435,0.00446724028449852,0.00452693242913571,-0.00697811262311832,-0.00698347652501952,-0.00219379185917579
"1269",0.00388083858176658,0.0157972723061393,0,0.0190887794122609,0.00463355649129649,0.000946430228110362,0.0052003073657152,0.00824950250529266,0.00778604193727372,0.00696219963645928
"1270",0.0110562632447802,0.0184857816222799,0.0120219644123587,0.0252245811635652,-0.0121047656041964,-0.00311964724567082,0.00638048177814188,0.0139391620854561,0.00685361993769473,0.000363970964420313
"1271",0.00527650280373249,0.0164218895391726,0.007559525957479,0.00876974878727577,-0.013753307441594,-0.00597542827593067,0.00633976954180882,0.0197253009046809,-0.00235151600180017,0.00436516390143638
"1272",0.0037272493338798,0.00255099678829795,0.0128616244248438,-0.00072448076155851,-0.0113254297620758,-0.00343470849416938,0.00476775612009339,0.00820600109046232,0.00527233590576648,-0.00724372798843753
"1273",-0.00257684961108962,0.00763348092686011,0.00423274770553239,0.00966658288562172,-0.00632625759665273,-0.00220166646866637,0.00305021541031025,0.00668637264833682,0.00672547018523906,0.0116745244053
"1274",-0.0011394952311472,-0.00280556996028791,-0.00948349572043894,0.00143612956347638,0.00180671677420952,0.00115125961425688,0.00557549114411371,-0.00779674940776742,-0.00704835113879987,0.00180315100471051
"1275",0.00836742448846306,0.00675260147655621,0.0127659679282304,0.011233338880541,-0.00240425513116493,0.0047914778232121,0.0127685297910285,0.0130964034424617,0.0272205612993197,0.00827933561250238
"1276",-0.00512956164043665,0.00251574433909907,-0.00210099216805193,-0.00401799619448417,0.0132565466769854,0.00534183113977593,0.00580629143676203,-0.00229785914877367,0.00510759530233873,0.00285608377297009
"1277",-0.000455018206593993,0.000557444237918592,0.0052632532292689,0.00522066146582922,0.00314303634693114,0.00303619200459537,0.00247414951039526,0.0051827602543002,0.0101631910046465,0.00356001051713029
"1278",-0.00341399596332503,-0.0153247233224688,-0.00628284769230603,-0.0144003209336655,0.0117714222799243,0.00340538775328914,-0.00872009578546562,-0.00773398889106869,-0.00556312951670035,-0.0102873049938557
"1279",-0.000380407898873947,0.00679140032529024,0.00632257144572312,0.00862282484149057,0.0115510460494301,0.00377086604606425,0.00514531946109775,0.00346390750536041,0.00761768141175789,-0.00250900001479271
"1280",0.00875724252656096,0.0207978852950701,0.0062828177608707,0.0220848504914937,-0.0114547208581642,-0.00347244229840815,0.00743061760583497,0.0161103256402333,0.00147658143614171,0.00323395006293814
"1281",0.00158522381272741,0.00220307166643319,0.00312169110409921,0.00278828474167203,-0.000419186916094771,0.00141659771005997,0.0021308409880556,-0.00141544136925964,0.00878747946198954,0.00250709217230694
"1282",0.0140185788818443,0.0189557575802115,0.00311209508278654,0.0166818315477226,-0.0214893044642432,-0.00791922372759513,0.0143931893509417,0.0144597897988905,-0.019935714353656,0.0117899484229973
"1283",-0.000668860696047102,-0.00620102888279539,-0.00310243999453497,-0.0084319251890741,0.00995114670354891,0.00275584210924351,-0.00483724106912531,-0.00614842794870052,-0.00274401099226917,0.00494350813762146
"1284",0.00252845697994442,0.00678240314709266,0.0103733043360581,0.00206843124951828,-0.0124011875296712,-0.00644457025798717,-0.000810159115714915,0.00337415739152735,0.0150735979514007,-0.000702731107745658
"1285",0.00296781358419618,0.00323359960476544,0.00410683885310559,0.00711011296411135,0.00077391816163952,0.00047709706208976,0.00064882266512134,0.00532534494775883,-0.00707128474492547,0.00457096435919468
"1286",0.00125753742723611,0.00268609609508763,-0.00306731207671773,-0.000455615688330302,-0.0074768776862385,-0.00228790599140805,-0.00729221039850925,0.00139386979413114,-0.00284864094955495,0.00525029928143272
"1287",-0.00738747940897311,-0.0192876688316977,-0.0123077892808063,-0.0221004492511967,0.0129883798903838,0.00563773853712912,-0.00832527733187216,-0.0153120596600197,-0.00523750136323065,-0.00940102202020787
"1288",0.0074424604321679,0.010106552940502,0.0103840465255056,0.0163091000906777,0.00128198186278161,-0.000665160473436566,0.0113578394408018,0.00706849571961343,0.00221368913613551,0.00246042320711748
"1289",-0.0012559580130278,-0.00892348685234834,-0.00308295699001493,-0.00825297211912523,0.00529281285916938,0.00209162148757769,-0.00992814337029224,-0.005614964612633,-0.00232821928028837,-0.000350626340403282
"1290",-0.00465991861958504,-0.00300156989484945,0.0164946802152952,0.00277388348947527,-0.00178307311748571,0.000759329204429893,-0.00493178008223838,0.00847018371171182,0.00592392310686707,0.00350749322354549
"1291",0.0110726386349054,0.0139573895308509,0.0101418227079026,0.0108345538690868,-0.00799646730925452,-0.00455107123540321,0.00826036421721477,0.00895828708079205,-0.000654339416725214,0.00454391175146429
"1292",0.00264642286182126,0.00431828637001086,0.00100427539548531,0.00182427382735995,-0.000257334030512868,-0.0010479503954639,0.00163854695719157,0.00721433594939103,-0.00386901190476185,-0.00173971176077381
"1293",0.000439968823371162,0.00134377017880194,-0.0010032678382802,-0.00409731215864462,-0.0110653264591911,-0.00362311280302807,-0.0124326711800307,-0.00688726862301692,0.0219300739074966,0.01568487205973
"1294",-0.00322415579966095,-0.00509912900205467,0.00301222350068131,0.00182874467617378,0.0125765103728954,0.0039236927677162,-0.00811627408297388,-0.00693459480263059,0.0112267451473103,0.00926559358588586
"1295",0.00441060471599464,0.00971109291296179,0.00600589670899199,-0.00182540647380303,0,0.00142980967053474,0.0116900592764189,0.00810024240405793,0.000462599740226777,0.00306014184494452
"1296",0.00219558786728391,0.00854927182604648,0.00199019388725796,0.0100570830643867,0.00651042295141369,0.000761199990912287,0.00280593856239997,0.0119146722982493,-0.00456599226526433,0.00610175144674652
"1297",0.00167992543769713,-0.00741733319065829,-0.00595841040437894,-0.00995694523905011,0.00885103452391678,0.0033287540111131,-0.00115223767574202,-0.0049288190870076,-0.00307727464616558,-0.00808621224280259
"1298",0.00291647080594748,0.00854072993586596,0.0159840881584372,0.0139430218137837,-0.00329025869523536,0.000473979265112723,-0.0075808320777585,0.00963154842209701,0.0104252069381223,-0.000339669258072273
"1299",-0.00392565507848097,-0.0108496231162235,-0.01769910235892,-0.00067619369808869,-0.00609379725752857,-0.0039793193446187,-0.00132843275010619,-0.00572393747541766,-0.0530290606654832,-0.0037377712839286
"1300",0.00518186850564084,0.0136436705902818,0.00600589670899199,0.00947419787344983,-0.00941431230648437,-0.00323965660814907,0.00532118894195999,0.00986862018593659,0.0141214200429116,0.0156890517662007
"1301",-0.00304968552534723,-0.011348716282093,-0.00995020149387005,-0.00245820621318515,0.00939225622160755,0.00401504913410244,-0.000330972141871055,-0.00488583439199708,-0.00162058098781237,-0.0100739096678047
"1302",-0.00407827294224505,-0.00400406263187525,-0.00603015629729353,-0.0172488010619912,-0.00793882741639695,-0.00199932908539802,0.00810721483351928,-0.00436457373686505,-0.00414814245877471,-0.00474902210510297
"1303",-0.0146251075093357,-0.0399358718534573,-0.00808901515020144,-0.0335083990579251,0.0121318502759116,0.00419778101409829,-0.0134581048635714,-0.0263014199585709,-0.0178086151937923,-0.0163598703524483
"1304",0.00697607015377066,0.0142379399910852,0.00611633038475667,0.0120284608526309,-0.00612079876973448,-0.00190031560827197,0.00432528389369047,0.0123803390090007,0.00571609107036442,0.00450444281824036
"1305",0.0099487963213285,0.0253232120062614,0.0172238673847416,0.0209741776403038,-0.0100078540823518,-0.00295067491089096,-0.00231882129548411,0.0216787079107188,0.0100836885019957,0.00827878144789507
"1306",0.00386733477180234,-0.00697958357612949,0.00398415267322916,-0.000456573629870505,0.0019870289023145,-0.000763851897620405,0.00464892490693769,-0.00516850103221667,0.00665540904317163,0.00273687664164446
"1307",0.0000727963430993128,0.00162197525448193,-0.00992061444010461,-0.0109615419479036,-0.000172135605228552,-0.000286642432413053,0.00694086805735794,0.000546634278952185,-0.00787353023579973,-0.00136470329624794
"1308",0.0180259257392428,0.0178134953339244,0.00901798576244683,0.0272457969919186,-0.0175936728798692,-0.00716743217861027,0.017889388211078,0.0177645240002331,-0.0167807831982463,0.00444138199630006
"1309",-0.00107106229663412,-0.00689441048015871,-0.0109237429460886,-0.0157340803960075,-0.0251951714595899,-0.0114540159466123,-0.00241854275076447,-0.00939835350402507,-0.0168206774463214,-0.00680273323384251
"1310",0.0057895992431749,0.0096128645517688,0.0080322803092685,0.00799269017253312,0.00153061695596124,-0.000292152133090084,-0.000646546956491911,0.00921653157667057,0.00946289987942417,0.000684922163946666
"1311",0.00138472051981275,0.00872766570095473,0.00597632865707842,-0.00113261570261325,0.00197843339354975,-0.000292237510902349,0.00598406073974234,0.00637943575600186,0.00136578716953339,0.0123204071609913
"1312",0.00391988354683726,0.00471944486275011,0.00297001594817781,-0.00385586282395733,-0.0119357524915539,-0.00613790235559619,0.00594861988269324,-0.00134293750382586,0.00179784869563826,-0.00169030813224702
"1313",-0.00291072109785762,-0.0117431069132015,-0.00987173393966745,-0.0173041093592842,0.00399666818726185,0.000490056742039391,-0.00239728343416923,-0.00995192692913449,-0.00903515710217606,-0.0121910687751201
"1314",-0.00163755008110933,-0.00580947476534233,-0.00498482184559867,0.00185352142576178,0.0113080384067226,0.00509474607612859,-0.00224299730755517,-0.00353153744722812,0.000499606554061893,-0.00239976354492633
"1315",-0.00720379273962701,-0.0114209233378697,0.0010019188574899,-0.0152638563559696,0.00321994355195976,0.0012676073896809,-0.0118816922711726,-0.0109047238658622,-0.00399475670705129,-0.00790370781297056
"1316",0.00323266243671427,0.00698531188942142,0,0.00751535924302993,0.00945224092112751,0.0036994158883692,0.00406235224791485,0.00303173007033819,0.0122829599173986,0.00969855199605174
"1317",0.0140353249946599,0.0170758018702168,0.00700701302177986,0.0174825894078388,-0.00512394333407751,-0.00116399476554274,0.0103334518783964,0.0129157212538107,0.0177675665063304,0.0044597718600301
"1318",-0.00310703493103659,-0.0115422799098185,0.00795232147503855,-0.00526925337193029,0.00719173448743704,0.00553599605234711,-0.000484778053033152,-0.00189922284625499,-0.00705589441809829,-0.00409837491775156
"1319",-0.00495847255419612,-0.0111466660022522,0.00197252914951429,-0.0168124320656575,-0.0014101221381404,-0.00173857852446835,-0.00226306348653948,-0.00679516438070105,-0.0105979536082469,-0.00960224010502808
"1320",-0.00170896692793565,-0.00778316631632747,-0.000984590245477923,-0.00117119804225141,0.0075032399760675,0.00415981880361582,0.000972071588676737,-0.00191585530905181,-0.00142403570751148,-0.0138504051469359
"1321",0.00413644614382846,0.0102786380250643,0.00295603412840184,0.00727007719549766,-0.0169102905198785,-0.00491366180283626,0.00841720580537331,0.00959706301809837,0.00520830856403953,0.0112359826673936
"1322",0.0073146518074525,0.01526104213012,0.000981925798251293,0.0137370399011216,0.00553989206568861,0.00239583244074715,0.00642064136534426,0.0103204591230508,0.00505802507580877,0.0128472255229006
"1323",-0.00408917577957413,-0.0208331199523238,-0.0127574223759721,-0.00574205249459347,-0.0173282184400344,-0.00735381915518285,-0.00462545086769861,-0.0129032445497825,-0.0187185648862335,-0.00445657267375199
"1324",-0.00991062854639302,-0.0258553808466193,-0.0228628993784543,-0.0180179963386635,0.0137457017422136,0.00506904829157828,-0.0100946179954406,-0.0152506879607111,-0.0167614736178715,-0.0154959387610798
"1325",-0.000500933005513904,-0.0091235356984406,0,0.00541056049379907,0.00722545602332092,0.00446095569190907,-0.00437043906835188,-0.00359497522133168,0.00699695280848123,0.0038475546290011
"1326",-0.0112306916821551,-0.00446429276275895,-0.00610365335203678,-0.0147402074816879,0.0233818034586544,0.0102350063628429,-0.00959191348497357,-0.00499600167714376,0.00669570471474579,-0.00452973397957102
"1327",-0.0167850166071795,-0.0252242011846093,-0.0122825952753916,-0.0194727598803673,0.011336582694585,0.00468309201122374,-0.019369528956263,-0.010878534039191,0.0108553118797552,-0.0133005924675427
"1328",0.00809432730878901,0.0169638636510199,0.0134715149610054,0.0108984435049655,-0.0119800496360988,-0.00390073630296595,0.0118848669298615,0.0118442665437899,-0.000186213525032453,0.0024831161464689
"1329",0.0130660140228473,0.0197907942929565,0.00511244984227521,0.0256347042028808,-0.00415703600896833,-0.0020051542302415,0.0142265219315336,0.013935490911869,0.0101197611545394,0.0130927143080344
"1330",-0.011888887363554,-0.0263377065619894,-0.0111900989960814,-0.0151833178873679,0.0161768144686203,0.00602865742923431,-0.00521934898949328,-0.00769643620268168,-0.011370565667558,-0.0101291689588564
"1331",-0.000656289018973744,0.0105351860140581,0.00205743835485372,-0.00498103494114444,-0.00145514696094229,-0.000285411068851715,0.0116413748393693,0.00332378952008616,-0.00242461290302975,-0.00988007454080853
"1332",0.0148124734906105,0.0208510320954141,0.00616037566989847,0.011442135251754,-0.000600259934083858,-0.00104625304442252,0.00858980998099135,0.0124241195463015,-0.00130878094751663,0.00463293958054045
"1333",-0.00337954946724028,-0.0080042599082143,-0.00204096371358864,-0.00471358482197859,0.00291637026862834,0.0020001396970375,-0.00530276484543368,0.00245416869749837,-0.00586584711388449,-0.00957784323772171
"1334",-0.0064209598435202,-0.00528701649577357,-0.00613485797365376,-0.0044991224533617,0.000940293953287208,0.00114065073230529,-0.000484810039651729,-0.00435246523375177,0.000753217007761098,0.000358161290763714
"1335",0.00167022760488322,0.0125876961489959,0.00205743835485372,0.00689826851879416,0.000171151103442346,0.0000943394779948648,0.0105060806782415,0.00928968796919172,0.000689958005580582,0.00393840047884164
"1336",-0.00840896807025659,-0.0223756981448031,-0.0112934986966602,-0.0191355557422509,0.0072606395621948,0.00199404023157523,-0.00927712211613974,-0.0143475875540182,-0.00294588203974666,-0.00178321596697351
"1337",0.00380131476522005,0.00734673755903215,0.00623041604219043,0.00216777064797347,-0.00703905327084919,-0.00255834398339849,0.0127542586131628,0.0120842704836495,0.00144587910906413,0
"1338",0.013691665663649,0.0165496612309435,0.00515993409217308,0.00913234926665507,-0.00512403494437597,-0.001235121838977,0.0109996309763838,0.0108551418662413,0.00200873819192582,0.00571639657127987
"1339",0.00696886078653636,0.00662274028938703,0.0051335632401619,0.00619189537426035,0.00600940453090226,0.00332947282497398,0.00425740011365017,0.00375842490947997,0.00883350485006607,0.00213140957556313
"1340",0.00164095687414822,0.00520815559642474,-0.00306441245845968,0.00142026711020282,0.00085321515438519,0.00104221832814511,0.00486708970001093,0.00401186560463862,0.00217354531561553,0.00319035098056442
"1341",-0.00370384727796058,-0.00627198290782327,-0.00204921153577609,-0.00212720941538291,0.000255474658932497,0.00085243365781329,-0.00140640793119118,-0.00372955712406198,0.00309827726179579,0.00388694552119162
"1342",0.00622008672787189,0.00768376885619015,-0.0102668036571638,0.0066315065734377,-0.00518602902851473,-0.00181973386004775,0.00876266129617997,0.00267370866547023,-0.00345934014518967,0
"1343",-0.00298428791176275,-0.0106208172023819,-0.00518669664601568,-0.0018821093452478,0.00704282303591586,0.00189920775575447,-0.00155132300131111,-0.00239968303283378,-0.00452523536029847,-0.0130235865097412
"1344",-0.00762527343497676,-0.00908338837902312,-0.00834194023427215,-0.00754350848355734,-0.00025598567489038,-0.0000950206163629064,-0.00341775483334772,-0.00908858768791865,-0.0100877703490323,-0.0110556673761554
"1345",-0.0161580572857083,-0.0172223712493785,-0.00736067828562625,-0.0175770850447534,0.00784822217047232,0.00398063831024698,-0.0076383656461696,-0.0129486644129603,0.00314524751119549,-0.017670375073744
"1346",0.000729731208219286,0.00819677941136865,0.0042370186930627,0.00362678236703151,0.000169486270126029,-0.000283627763522198,0.00565505542108435,0.0081992483002169,-0.00244559476738193,-0.00220261312828607
"1347",-0.00401157591994172,-0.013456814466684,-0.00843864604757605,-0.0158999163236693,0.00533165108316225,0.00226619105963977,-0.000937234167778578,-0.0103011302766454,-0.0193613399627692,-0.00367920130409782
"1348",-0.00593179238378694,-0.0147769491594799,-0.00851064528548673,-0.0129744034940382,0.000673436749148992,0.000848264721812431,-0.00234501644961804,-0.0106819662951885,-0.00980768589743597,-0.00775473278825167
"1349",0.00206300458874153,0.00519202101928529,0.00429178770743599,0.00421630572552312,-0.00294456599351056,-0.00141184684296181,-0.000940382704538889,-0.00027674606298167,0.00194214409307869,0.000372080552337062
"1350",-0.00301446992779941,-0.00487802807909676,-0.0106838312236726,-0.0128425929562263,0.00826895914179215,0.00329894858237667,0.00423521236453106,-0.00498493350747164,-0.00781809115931786,-0.0074404513480204
"1351",-0.0110610908381678,-0.020472988786025,-0.0107990846655361,-0.0227669614580341,0.0139744235159915,0.00441568050958097,-0.0121835532702826,-0.0125244855554021,-0.0145219850810365,-0.0131184545155544
"1352",-0.00574157784951423,-0.0156019968514644,-0.0131004485367051,-0.00870484369422664,0.00404405871842473,0.000280376854818076,-0.00490189628046056,-0.00930053757599858,-0.0105068193946103,0.00189894864774565
"1353",-0.00382489959625232,-0.00687799113216725,-0.011061830566068,-0.0142044469706305,0.00287734329066902,0.000748241346059997,-0.0122357013020432,-0.00825067382790357,-0.0018698944213339,-0.0011372096858524
"1354",-0.0148310850114772,-0.0165613693439631,0.00894871288293064,-0.0136232375431488,0.0177029202033925,0.00373743791519243,-0.0276707236750848,-0.0117610648944485,0.0223470884756483,-0.00227693068930646
"1355",-0.00855867438097702,-0.00275567866019411,-0.0144126161269644,-0.00956176816748833,0.000241799098012363,-0.000651538224474946,-0.0102581306823021,-0.0072569485552938,0.0114528793562916,-0.000760813374248825
"1356",0.017188189301536,0.0239485165530484,0.0101231642323738,0.0238670579421942,-0.00209357438325319,-0.00260860294708698,0.0205616938989093,0.0236839152499446,0.000646981546807091,0.0133231960579028
"1357",0.00174265914978888,-0.00329834617630265,-0.00111304617312902,-0.010476458037591,-0.0111341936450928,-0.00214739583136125,0.00212925071799064,-0.00628373022770179,-0.0166181189764546,-0.0142750178179645
"1358",0.000530021208825504,-0.0105292953172792,-0.00780373339329399,-0.00688226521061974,0.00693539387734576,0.00262021199576945,0.00424969896672112,-0.00546148757362896,-0.003024769818191,-0.0110518353072266
"1359",0.00196561606093804,-0.00638505493460484,-0.00449454621835654,-0.00506371966926211,-0.0038084853299154,-0.00214680750480656,0.00309274874619581,-0.000866892209536174,-0.00138498223799577,0.000385351197087491
"1360",-0.00324481372140173,-0.00152996047320086,-0.0056431850076174,-0.00482184967713783,0.00374199672464171,0.00290001733159517,-0.00292073922175218,0,0.00838774827586697,0.00346682482868865
"1361",0.0121120080826194,0.00950042400677642,0.0124858541510124,0.0282634283854628,-0.00307954853710213,-0.000840043115964861,0.0136695315569695,0.0138846658243947,-0.0108723413420644,-0.00422251234308701
"1362",-0.0145101037815978,-0.0258045796003582,-0.0134529892355577,-0.0172773546857622,0.0253615404567937,0.00952307924133811,-0.0232781736153163,-0.019971349164595,0.00589325901487858,-0.0185043039401039
"1363",-0.00220093251344133,0.00124665647630784,0.0102272813646407,0.00426223703029049,0.0115743435488858,0.00388446894408578,0.00624582378530669,0.00378454149904472,-0.00190908427597691,-0.00864096828130689
"1364",-0.0251767066416628,-0.0211641306544933,-0.0269967444515005,-0.026790404727279,0.0237406056264688,0.00859039611285928,-0.0253184399294298,-0.0179810911268716,0.0387811976909775,-0.0206023441985491
"1365",-0.000468151960336338,0.00699522059095647,0.0115607708119039,0.0043607840710711,-0.00790159699544457,-0.0057632268888681,-0.00703864081330341,0.00383912265542175,-0.00114281269841265,0.00566352009082416
"1366",0.0075721742017969,0.00315754683418334,0.0125713416558173,0.00271368480697509,-0.0133766408724788,-0.0033128729870624,0.0197467223153078,0.00617834589207455,-0.00114421556058042,-0.00362030687199211
"1367",0.0224682654487434,0.0336794513494432,0.0158013374330723,0.0292286345838344,-0.0199842313637827,-0.00655467418801037,0.0213507660452286,0.0362569229353018,0.00044551355762712,0.0185708895967318
"1368",0.000606364433778817,0.00182714110277993,-0.00666648266702763,0.00604780785148296,0.00151947246843664,0.0024160939762381,-0.00486149927334711,-0.00423207961248973,-0.0172381329389546,-0.00673799981177947
"1369",0.00795133360162836,0,-0.00894871288293064,-0.00862509784390231,-0.00023923906034784,0.000741692407574712,0.0125386445793454,-0.00510062983160531,0.00148864724919084,0.0031922947283809
"1370",-0.0126968718100294,-0.011246266834669,-0.00451448348121042,-0.0145003236724489,0.00455222733770033,0.00268629518656516,-0.0196206023114716,-0.0150954087703612,0.00407164102815605,-0.0182974890606896
"1371",0.0114906328954589,0.0190594593902209,0.0113378772994333,0.0208666810729969,-0.00914374791822414,-0.00535837987761489,0.00935045050030947,0.0118567462956414,0.00708036813156299,0.00486217012124057
"1372",-0.00639501995993974,-0.00904984537704057,-0.00560554570408034,-0.0036688750811168,0.00986995801020618,0.00529433950284686,-0.00471331707167355,-0.00600235162869778,0.00421825367807882,-0.00766118603546284
"1373",0.0106005302593293,0.00700167977519262,0.00789190629084757,0.00710157659718247,-0.00127163276523579,-0.0026791088271011,0.0135532352358678,0.0112133928974325,0.00400970608483031,0.0117837915331112
"1374",0.0102272882630998,0.0157192566949607,0.0145414625956386,0.0182814693322879,0.00556892286070543,0.00463207026140644,0.00628353165532669,0.012037773223049,0.000570497622820909,-0.00160644505840102
"1375",0.00193801319252551,-0.00922615746370403,0.00220523084045565,0.00205200265730321,0.00537999755349428,-0.000276566414039725,0.00784486279502583,0.000855107845812331,0.000570178676385646,0.000804494238004771
"1376",0.00967276121326988,0.0231301537919149,0.00550017581518847,0.016124690208027,-0.0130626342290288,-0.00341306634100891,0.00466380267874267,0.0170991966206899,-0.00487550835261552,0.00844052334810597
"1377",-0.00162120225033602,0.00703779031734619,0.0087528685381546,-0.00327437954167742,0.00494348785626975,-0.00203629602712618,-0.00127635159711925,0.00196109827036373,-0.00757192014324448,-0.0163411536663084
"1378",-0.0224387816754482,-0.027594626358544,-0.0144548687341233,-0.0366221755220169,0.00531528957062588,0.00213289584109289,-0.0156522924651221,-0.0209734768547958,-0.0253253636896495,-0.0214749183216139
"1379",0.00770159403802562,0.0111042815365778,0.00666705946529822,0.00318559056915935,-0.0133372561508666,-0.00434978111669704,0.000811039027299953,0.00942637009240888,0.00407837773770869,0.00993788052228783
"1380",-0.0160345425608525,-0.0265405275210185,-0.0154526826669585,-0.0185235404167606,0.0145576075333118,0.00548414324262492,-0.00551223427677527,-0.0116014963177707,0.00733750004807066,0.0102500893865118
"1381",0.00502569010703002,0.00626757601820693,0.011210891140395,0.00862765357491324,-0.00394222304581704,-0.00221814111307439,0.00440183637693314,0.00973350591015532,-0.00741415216617314,0.00689934024072114
"1382",0.00901674334026481,0.00840874066463826,0.0077606987977985,0.00641542995114963,0.00158326652286389,0.00138945254826028,0.00633004006540361,0.0110574372935379,0.00137601236325557,0.00564301657149979
"1383",-0.00285375964277446,-0.00154420809619982,0.0143012009511729,-0.00478083021717013,0.00245020227852599,0.00323838494345541,0.00838726217286201,0.00168291236512275,-0.0116469212635357,-0.0108217008893704
"1384",0.0249268998917598,0.0423754798338514,0.0206071347121577,0.0443022353486329,-0.0130077822471679,-0.00461097747203687,0.0227125003363449,0.0296750216100696,0.0274081358343303,0.0433548923793641
"1385",0.00301256822913931,0.00919871841714848,-0.00318799954653148,0,0.0103175834839153,0.00463901614702666,0.0106351823061384,0.0103317404693373,-0.000644410069663981,-0.00194172110753565
"1386",0.00659259082590036,0.00793890523750163,0.012793204130586,0.0199335399491622,-0.00768484294540317,-0.00249350649015356,0.00557097038602339,0.00430574058887601,0.0152815208016381,0.0280155820911756
"1387",-0.00451176881493864,-0.0239204927688609,-0.0126316054239011,-0.0105238416236325,0.00510966740758767,0.00268535246351109,-0.00461667213523487,-0.00911037324150166,-0.0113045466840351,0.00378503751243242
"1388",-0.0095036939070785,-0.0128511509439094,-0.00426432088874329,-0.0182323475688335,0.00929398796916669,0.00350893900115867,0.00139125158320952,-0.00432674022920509,-0.0126540730252988,-0.023001542465737
"1389",-0.00125499230482107,-0.000605618582688261,-0.00535351696406972,-0.00361128897087049,0.00881478403972213,0.00276046755119719,0.00200741870584742,-0.000814736796939663,0.00214680882813312,0.0177537984865639
"1390",-0.00871988474710117,-0.00424114166440948,-0.0107643884535809,-0.0111310062677402,0.00202835549201907,0.000459030506535063,-0.0118647320370618,-0.0103289735121278,-0.0122695344448635,-0.0128934580304473
"1391",0.000149110384929152,0.00365090517720867,0.00217658153901357,0.00523549927768552,0.00124567589208291,-0.000917479533711907,0.00155958350982432,0.0107115671484312,0.00552094007969539,0.0111409573662571
"1392",-0.00484516292805648,-0.0103064071285452,-0.0152007362147177,-0.0166664026987098,0.00707624991755651,0.00229555389229508,0.00435934230577617,-0.00625035190354084,-0.00261460871251018,0.00227960414753747
"1393",0.0167776613087314,0.0159265537462945,0.0099227012811367,0.0193325497753987,-0.00262557753326809,-0.000825127208756049,0.0108509473309546,0.0150398692909448,0.0101579595034524,0.0121305097542026
"1394",-0.00235723712854152,0.00060310023595278,-0.00436695515953089,-0.00233846179574271,0.00464523305806308,0.00220068986768962,0.00383356356635089,0,0.000454184510537026,0.012359496595415
"1395",0.00686690270972878,0.00421791416558981,-0.00438598492718734,0.0132811523119556,-0.00785988368114909,-0.00256116248800831,0.00840213653459965,0.00942874649218162,-0.00479868988009313,0.00110978658825989
"1396",0.00740738057689527,0.00690091481115518,0.00330414359793307,-0.00257005947460953,0.00054361498447042,0.00100882132232383,-0.00772596818474192,0.00400338786528254,-0.00273667816031353,0.00886924934503464
"1397",0.00262044854485843,0.00953504338807365,0.00768393658217947,0.0092761455829582,-0.00256174085380534,-0.00146574727703663,-0.00839708655111671,0.00318964444954251,0.00215617114362288,0.0120879356194799
"1398",-0.00914824955429572,-0.0242029794191546,-0.0239651375135557,-0.014807337861561,0.0122186713173462,0.00394501755480237,-0.00338717778595954,-0.0116584364486747,0.00189068320867491,0
"1399",-0.0101123592594033,-0.0229885774597075,-0.0133929783150454,-0.0261725559046556,0.00561278427846079,0.00164534545724138,-0.00602518209351566,-0.0131370545777925,-0.00416476220686868,-0.0209916867428366
"1400",-0.00858640775184272,-0.0145510979697042,-0.00904978201596318,-0.00425759509840207,0.00787537960468909,0.00191604635527609,-0.00404103840430636,-0.00869298540770469,0.00320201923284325,-0.0059150056241617
"1401",0.000223813794808958,0.00691158254727897,0,0.00481040512161268,0.00257907403077628,0.000545825161954561,-0.000155929981033975,0.0112358263140073,0.0140046504949283,0.00743779921520837
"1402",0.0164973403321305,0.0390016899124044,0.0148401437988483,0.0226063081143553,-0.0091557074732278,-0.00309443155610356,0.00811619827772092,0.0181570767953865,0.00706626847904257,0.00184567420582926
"1403",0.0184330112961477,0.0252252411879983,0.0179977675479173,0.028088245417631,-0.0188617875148768,-0.0072124033354134,0.0113019619037225,0.0159703522140611,0.00491158372363132,0.0103168479898337
"1404",0,0.000292964029978249,-0.00552503523476566,-0.00581846982379308,0.00747178584780639,0.00321869223874205,0.00275582163692012,-0.00314412863171176,-0.000698235399820168,0.00583515216558039
"1405",-0.0069947536054189,-0.00732063789251258,-0.00111091967508115,-0.00458004915629984,0.00200868732576143,0.00174148096316684,-0.00106888027527652,-0.00210221033756652,-0.00597083174614632,-0.0119652153326775
"1406",-0.000871460608794061,0.00147496922031043,-0.00333690646452045,0.00178930862237592,-0.00499873886894453,-0.00364767314392977,-0.00290383924959992,0.00237030402181282,-0.0086267873785294,0.00146794543273732
"1407",-0.00690466014247604,-0.0191459177228694,-0.00446436823550822,-0.0117374156466469,0.00566832369224146,0.00239218357818705,0.00107274576139305,-0.00236469896634262,-0.00651021017474662,-0.00842810650609738
"1408",0.019833347826627,0.0441440969998523,0.011210891140395,0.030983552837998,-0.0161375781172819,-0.00523035009803374,0.00734983928856625,0.0265995366987142,0.00921298873635923,0.0169993723911357
"1409",0.00193744133765583,0.00603958562463003,0.00997770501485107,0.00626139044116503,0.000392201733881992,0.000645450810315529,-0.00288811402378419,-0.00307804324665018,0.00482160067846471,0.00581391130596076
"1410",0.00501390069595087,0.00857633092479038,0.0120747042103964,0.00273730940975625,-0.0128657759697636,-0.00525461981577502,-0.0103657506725938,0.00386010849609764,-0.000127984642457113,0.00758667603917651
"1411",0.00121134020077274,0.000283568416735713,-0.00216937570969222,0.00198538939713844,-0.00532462031237957,-0.00139003389828973,-0.00600746503218963,-0.00589605772402702,0.00127973509905122,0.00286844636302375
"1412",0.000854090352912174,-0.00113359788673717,0.00217409213235475,0.00421134020089764,-0.000719242903936324,-0.000741966038616648,-0.0029444231163599,-0.00567298886288792,0.00325926005263955,0.00822316790061595
"1413",0.00163590855880047,0.000567513120482754,0.00108447290707736,0.0046867029717641,0.0050373941199382,0.00287886790767122,0.00217598747934078,0.00207452551565557,0.00121019169341396,-0.00531922193021361
"1414",-0.000497117900488786,-0.00255177573776855,-0.00216681091419235,-0.00883895659873601,-0.00167068934773262,-0.000648036539641517,-0.00031011438605788,-0.000776561133836062,-0.00757086176992006,-0.00784314027661215
"1415",0.000142020589903868,0.00454803669883597,-0.00108586568016122,-0.000247198318910735,-0.0135468064764358,-0.00491156991896435,-0.000465389424708307,0.000777164649697459,-0.00551317374468951,0.00107795869947758
"1416",0.00113658947001216,-0.00226381128630848,-0.00543489182146795,-0.00148698673327341,-0.0140561153091117,-0.00502842836967676,0.00279372076717643,0.000776521205760883,0.00322310309988061,0.00861456835818042
"1417",0.00737850748252855,0.0116280071516934,0.0131150623999152,0.00918104359468219,-0.0085210645423095,-0.00243337410616917,0.00727433448140147,0.00517166083863208,0.0059756664532653,0.00391453712345635
"1418",0.00133828373732214,0.000841123565295643,0.00755115872239687,-0.00491744724374987,0.00487563206469521,0.00121993861616465,-0.000460726878704576,-0.00154349586591818,0.00102199158178307,0.00141799052216385
"1419",0.0000702065777147265,-0.00224094771520023,-0.00214138253578322,-0.00049431514196896,0.0020558027539328,0.000562300511121494,-0.00076879427355081,-0.00206124215967896,0.00344559722150595,0.00460174330616092
"1420",-0.00302439945859179,0.008422305322211,0,-0.0014832108025602,0.00443196158536585,0.000842846061281932,0,0.00180732713605081,0.00998351169984457,0.00916132853008333
"1421",0.000423851387851393,-0.0025054599977643,-0.00107292819297444,0.000495177055165774,0.0165042618204807,0.00776594703672928,-0.0009230670490048,0.00180398707068363,0.0107661712426346,0.00523746664346136
"1422",-0.00817957068676456,-0.00586118751672715,0,-0.00915613907732016,0.00417993892275659,0.00176463612999767,-0.00261783211480637,-0.00565957745595036,0.00840915696314992,-0.00486276892515303
"1423",0.00604272233367631,-0.00364948197816028,-0.00107420224426902,0.000249797086041337,-0.000960948709704423,-0.000463595657057225,0.00385983665697576,0.00129365408939863,0.000494175060190116,-0.00453753155768599
"1424",0.000211766929127943,0.00338095906495361,-0.00322561554651879,-0.0102372024702612,0.00584907829437253,0.00259641016768941,0.00215300088559855,-0.00310098972939921,-0.0037661295069078,-0.00455828677532077
"1425",-0.000989002518853255,0.000561916240042981,-0.00863039306797853,-0.00201803440458059,0.00238987506269028,0.000370285564455397,0.00399018455674094,0.000518592592172018,0.00173523796643993,0.00070453633450196
"1426",0.000778049918792378,-0.00336830587143377,0.00326481069436824,-0.00480292341248401,-0.0043705666396241,-0.000647673860630804,0.000306051859785939,0.00259069966917269,-0.00649593545221427,0.00175991964506861
"1427",-0.00720803080304999,-0.0121088327321672,-0.0184383117252995,-0.0116841998839667,0.0051880970147864,0.00185061854291657,-0.00106979817313435,-0.0108526069303263,-0.000435842840422085,0.0010540966616186
"1428",0.00476871588666627,0.00940700725541599,0.00110518849207453,0.00950923526080838,0.0141332255028084,0.00646380948659897,0.00397736526176873,0.00783666545070827,0.0230500679529013,0.0105300477460186
"1429",-0.000920491816817748,-0.000564983937814456,-0.0132450896093098,-0.00560075035336616,-0.00100424258196186,-0.00228765919130203,0.00502820651381586,-0.00596145538963988,0.00158321153584695,0.000347338084005111
"1430",-0.000850560830947034,0.000565303325113176,-0.0123043433332823,-0.00512034843900078,-0.00471241848441739,-0.000368172115287391,-0.000606537972958954,0.00286835909736571,-0.00103354817688583,-0.00486111622344032
"1431",0.0202962696653999,0.0293700566773782,0.0135899657457361,0.0221307335644161,-0.0166506973191752,-0.00681724486398827,0.0078884229762064,0.0176803391220797,0.00352991909841038,-0.000348877680432791
"1432",0.0038950085575038,0.0145406374742061,0.0134080078824823,0.0231621575641328,-0.00465490169521587,0.00129841004691822,0.001806325363918,0.0107308455046315,0.0215295228426802,0.0111692034417417
"1433",-0.00568138410792329,-0.00919431793247627,0,-0.0127951409623217,0.0024188625335384,0.000463191100611438,-0.00646028977013446,-0.01238632517752,-0.00682741027276867,0.00138079096165633
"1434",0.00278738792369349,0.0136461750741059,0.0044100374338607,0.0119638417752514,-0.00627328719464848,-0.0018517345574709,0.00393132676317975,0.0104942239969295,0.00364636873408197,0.00206822407648244
"1435",0.00333534354917453,0.00376972550945665,0.0109769190705422,0.00443342566831717,-0.012464564734786,-0.00491638969012709,0.00376565189474465,0.00531929257058739,0.000119142350892609,0.00515995919531664
"1436",0.0152360842716768,0.0160943862774763,0.0162865096743765,0.0269741357191369,-0.00393443326848641,0.00288991729032495,0.0121549254156414,0.0191481166375407,0.0201881850903787,0.00684463933566049
"1437",0.00443481310516058,0.0116156633217896,0.0106838850993929,0.0117001139752484,-0.0265771011859764,-0.00938859853996288,0.00518929120184053,0.00321406405807756,0.00286034093585119,0.0105370807807292
"1438",-0.00339623467777717,-0.00443650052695632,-0.00951365716046149,-0.0108570145082556,0.0120024756669388,0.00206457134714211,-0.00472011836305453,-0.00936428986245597,-0.00814906272149485,-0.02758157108499
"1439",-0.000817584177888908,-0.00786366415765105,0.00213443569857241,0.000477641477642843,0.00501195808274013,0.00252811590938351,-0.00859496094019807,-0.00273631916216699,0.00774652022581646,-0.00726389441688557
"1440",0.000545360076979584,0.00660494887486784,0.00212973883171541,0,0.00656594995825133,0.00233493701690746,-0.00463393750312935,0.000498828683903829,0.000116491962983467,-0.0146341610358031
"1441",0.0000685978993548719,-0.00839878308349029,-0.0106268456760304,-0.00596250394011422,0.0024770299093404,0.00055975481094217,-0.0117133050020268,-0.00299178758538921,-0.0015721671837613,0.005657667601356
"1442",-0.000418252162818766,0.00158809554368733,0.00537043343166488,0.00239914280275033,0.00115314471912398,0.00214169238111639,-0.000303991079744992,-0.00317904418026893,0.00285767771121659,0.0066807125953503
"1443",-0.00150801779365661,-0.00369995611878937,-0.00213659553463419,-0.000957405590012672,0.00781582378350265,0.0022309119025099,-0.0010641070232339,0.000759627789736594,-0.00529195140123473,-0.0104784481678606
"1444",-0.0106421373584905,-0.00822266197498789,0,-0.0148537244782269,0.009877543876184,0.00370936077242279,-0.0146786421968976,-0.00758749537509373,-0.00163694238578882,0.0010589336079363
"1445",-0.00562106594201972,-0.013104949726814,-0.0107067308050809,-0.00462048179943619,0.0107507228741086,0.00415702268298856,-0.000933729451598642,0.0033131095878276,-0.00562163130241533,-0.00705219856480976
"1446",0.00942140428374771,0.0121951037732257,0.0119048538258537,0.0158805963797968,-0.00711789987203826,-0.00211624916289432,0.00545310186884618,0.0099058082839476,0.0148989931676462,0.0124289901219379
"1447",-0.00463210384776624,-0.0222221523091745,-0.0192514672800239,-0.00601249526763403,0.000564147664566361,0,-0.00232429129698863,-0.0128269745680026,-0.00261110021146815,0.00596284678055925
"1448",0.00263965089030482,0.00930992233904204,-0.0032714675916431,0.0099200396774104,0.00371106420470557,0.00185613090188097,-0.00714506965920081,0.000764270105686027,0.00232703474505236,0.0013946092478001
"1449",0.00103884292269707,0.00623965497863654,-0.00437617037420812,0.00143759803173804,-0.00136624922481654,-0.00064551365604204,0.00844796739198239,0.00229152648684305,-0.00110271639514203,-0.00522287761086537
"1450",0.00408319068110341,-0.00269615590842731,-0.0043955920876606,-0.00669860341049866,0.000321914255806854,0.00101441961618387,0.00294769792019567,0.00101592058170197,0.00180126664260527,-0.0171508047357199
"1451",0.00716783428425116,0.0121655016771489,0.0121409962139836,0.0103564591614058,-0.0124709061366969,-0.00396086978614929,-0.00371231152789209,0.00888086544825351,0.00696013556150743,0.0217237170535389
"1452",0.0000686201597974723,0.002136901315132,0,0,-0.0129544172568382,-0.00453140815922071,0.00434711252722897,-0.000754428372629623,-0.00570247102296839,-0.00522833851815707
"1453",-0.00342120074632946,-0.0079961010686278,-0.00545257977453695,-0.00882001380618069,0.0084190200693528,0.00325112127434934,-0.00417379946922924,-0.00402713050699455,-0.00330200449837803,-0.00280311720481063
"1454",-0.00988772721425246,-0.016388754358613,-0.0164472649766633,-0.00745528355153635,-0.00180041904827444,-0.00203713784806769,-0.00434658410343525,-0.00657061032358741,-0.00616098797743125,0.00737878512213519
"1455",-0.00638003489386241,-0.00273150537544464,-0.00780373840625048,-0.00605777149905518,0.00705225735829118,0.00241277759798275,0.00124741640420445,-0.000254251110860748,-0.000877296892294877,-0.00174399536590708
"1456",0.000558546816228356,0.00986012698098993,0.0056178988944251,0.00926372146483634,0.00692128777296297,0.000925630547964129,0.000155481706220373,0.00610684694241126,0.0028097109063383,0.0115304929006563
"1457",-0.00327831902565578,-0.000270966710356424,0.00111747370341697,-0.00313994216616531,0.0025065391267185,0.0000924002222411069,-0.0043588987514549,0.00126432473700544,-0.00735471018279843,-0.0138169849865292
"1458",0.00832758359108254,0.00922387760651477,0.00669647335858792,0.00581516131856774,-0.00225851966138568,0.000277153604169245,0.00672381491561813,0.0101036412822832,-0.0100552276849962,-0.00490368285955811
"1459",0.010133185277444,0.0185484864181977,0.0144120627134694,0.0103589536747304,-0.0138249400724263,-0.00471469141245673,0.00465989246768039,0.00975234513770418,0.00635575860923931,0.000704040312520915
"1460",0.00453540799223773,0.010293016004628,0.00546459128394483,0.00786847631653509,-0.00926361031137735,-0.00631602259129427,0.0015460651632988,0.00990585874475691,0.000708269398043582,0.000351663888966014
"1461",-0.00259925901517122,-0.00548592901594769,0.00652147628389144,-0.00283911694883254,-0.0061236957857228,-0.00177596189180829,0.00941627105336518,-0.00662096300178028,-0.00442373499449178,-0.000351540264949435
"1462",-0.0166645992099289,-0.0133964765822788,-0.0129586583994451,-0.0154212575230449,0.0135711619880177,0.00421380152698614,-0.00932843200906497,-0.00987407105480886,-0.0107825823536826,-0.0151249139891453
"1463",0.000139625660130038,0.00559099152410103,0.0142233435938965,0.00963882449371001,-0.00640694906350503,-0.00335682670744997,-0.0035502469842098,0.00772850930456581,0.00365335686857904,-0.00464283041474622
"1464",-0.0138763788408559,-0.0238284386572624,-0.0204964734535746,-0.0205251524719562,0.0143021479322123,0.00477135527317296,-0.0100701702651693,-0.0113802785143957,-0.0128297468333961,-0.0121995151716672
"1465",-0.0028287516661083,-0.00135581678934427,0.00220294948033084,0.000974755226418322,-0.00986261240733466,-0.00214197779099556,0.000626092834170588,0.00400418139752623,-0.00344551788743641,-0.00290588105193434
"1466",0.00290769165710469,0.00624667091436137,0.00769203725942846,0.0109541294138606,-0.00510365463357776,-0.00363927163175715,-0.00437898294971895,0.00822516052974898,0.00703629135608219,0.00255005608008707
"1467",-0.000565844635537993,-0.000270021314577762,-0.00545257977453695,-0.00770529435770939,0.0147281133395578,0.00636899788994993,-0.00581214610202074,-0.000494284633097086,-0.000542169605055598,0.00218020271517072
"1468",0,0.00242993698565908,-0.0065786514337316,-0.00145585722038855,0.0058709439728899,0.00409509660530682,0.0112182919498931,0.00766733757462146,0.00542402843348522,-0.000725227892248381
"1469",0.0104705269775729,0.0115806137942129,0.00993340315633473,0.016282015999219,-0.00818720852835941,-0.00199548560299534,0.00109341477050329,0.0108006098938316,-0.00455550554989503,0.00181427353995822
"1470",-0.00889150640215108,-0.0122471699576354,-0.00765022358198131,-0.00526066479171383,-0.000735995840636994,0.000837218976179166,0.00671162263861769,-0.0111707254471298,-0.0208948085369804,-0.017022771955908
"1471",0.00204842088034707,-0.00377352044098622,0,0.00480762639623689,0.00564360969879862,0.00241543260140875,-0.00744195241906098,-0.000982239660393569,0.00387447710180266,0.00847457402154794
"1472",0.00782534874746954,0.0113638135457501,0.00220294948033084,0.00789494333442531,-0.00943450269261792,-0.00454193749054255,0.00218683947073228,0.00958692930735849,0.0188078605356334,0.0179027562684033
"1473",-0.0226637518916307,-0.0160515974948082,-0.0120880960232966,-0.0163782493985535,0.0181456676714402,0.00838075357060442,-0.00498760710987423,-0.0126613766373163,0.00114252553561278,-0.0186646826118815
"1474",-0.0120239799680589,-0.0108753191148472,-0.0044494080714218,-0.0125481049282979,0.0148388515141464,0.00443278220936438,-0.0101816022223421,-0.00838483182877592,0.00900954985255731,0.0014629624526632
"1475",0.000869228776379627,-0.00329872876907877,0,0.00195514057681967,0.00111266290018963,0.0000914881437392712,-0.00332346216671953,-0.00174079757925893,-0.00101195306232649,0.00803510311144295
"1476",0.000796285637732819,0.00193084827904655,-0.0100559980035667,0.00365841417945645,0.00166681518587342,0.000643584863952995,-0.00158794737106993,0.00024895576675088,-0.00220480267290191,-0.00471015522293972
"1477",-0.00347165724285325,-0.00330337151103233,0.00112876125801464,-0.0089915992700238,0.00332814104143742,0.00119451654430058,-0.00318041168478356,-0.00423397495248545,-0.00209012246205054,-0.00182014263204167
"1478",-0.0134988929863802,-0.00938924979523714,-0.0124012892897808,-0.0154484565398149,0.000947944060496253,0.00027497721189218,-0.0194638439188093,-0.0120058856355381,0.000239335718515754,0.00291761361802267
"1479",-0.00169187262473025,-0.0011152330074119,0.0159817902796966,0.0034867226457469,-0.00197270049195186,-0.000458442097421186,-0.00439295455189415,0.00759494866578736,-0.00628217665598985,-0.00400002006035627
"1480",0.00493732965233717,-0.00558193714836175,0.0179776709172168,0.00297840714291464,-0.000869788708135033,0.000642277021456028,0.0114396088843174,-0.00175873012116268,-0.00126432057954895,0.00438110108307055
"1481",0.0202392752510239,0.0224529048528759,0.0143483080296829,0.0175699533921243,-0.00561823519903615,-0.00201743800077381,0.00937148816157696,0.0148505513167105,0.0119965634194428,0.0189023340870691
"1482",0.000430851230274421,0.00329385800535054,-0.00217608862579644,-0.00194563109925072,-0.0100272228087673,-0.00413600937339043,0.00624277387518513,-0.00248052829848355,-0.00285933171082775,-0.00677854216455243
"1483",0.00186793361201487,0.00355675939046352,0.00109072589988357,-0.00194910681554528,-0.000562884043231127,-0.00147672529106235,-0.000636515493969592,0.00124317722001122,0.00101558636128574,0.00431032299677248
"1484",0.0136250271922393,0.0239913174130533,0.0119822911911749,0.0163573384072178,-0.00096472966354022,-0.000554251065958855,0.00811888597000388,0.0144029579269298,0.0122344415401581,0.00357656282013474
"1485",-0.00212228092192679,-0.00212997443617979,0,0,0.00474982138196522,0.00166466073535965,0.00142095261260611,-0.0019584144722552,-0.00106130534130477,-0.0014254239409307
"1486",-0.0051044017525298,-0.00586968235868734,-0.00538202661177845,-0.00840729775819682,0.00392629902904962,0.00230804090074965,-0.00536117726441498,-0.00220755362385805,-0.00424946012952976,-0.00142760560061006
"1487",0.00805219357580333,0.00939328939084705,0.00108224829676362,0.00557157421120547,-0.0014367797636764,0.00128925349990405,-0.00174357256254298,0.0054077049006489,-0.0128030579715404,-0.00321664961115631
"1488",0.00466547178053811,0.00904010836802649,0.011891830710502,0.00722721808229765,0.000159845910218559,0.00101201850152965,0.00651100203699539,0.00831315541169042,0.00378258774333373,0.00681249553246777
"1489",0.000211239981745326,0.000790490945340894,-0.00320493867326233,-0.000478359232643055,-0.00271719950838889,-0.000183616061264047,0.0039445588269027,0.00193996868700186,-0.00675912218754549,0.000712314306763551
"1490",-0.00492437256667833,0.00368621950108072,-0.00428747662464657,-0.00047858816971269,0.000923373600630217,-0.000395810527934026,0.00282873851181997,0.000484210407111663,0.000481794631464139,0.00249106907856311
"1491",-0.00141373208268369,0.00524680921966403,0.00107651503399975,0.00287279064669166,0.0057759514274407,0.00174905951652615,-0.00125361465525475,0.0021768935461659,-0.0102931857493174,-0.00887467772603245
"1492",0.00176982465890774,0.00182678857783958,0,0.0107423169526111,-0.000478312790886171,0.000827221501987996,-0.00266762276758536,-0.000482703327611578,-0.00182461381613697,-0.00107455759836994
"1493",0.00339208750459652,-0.000260661392872841,0.00537645210845117,0.00755810946043045,0.00215417549659369,0.000550961442270514,0.00881041045364839,-0.000241652858283703,0.00231540952703546,-0.00896381185338879
"1494",0.00302885330451486,-0.00286600351406496,0.00320848704034482,0.00304722885761,-0.00923653371769484,-0.00284492857089991,0.004055074527481,0.009420201743217,0.00401218237082057,-0.00108533151390944
"1495",0.000421438339263336,0.00130654449473377,-0.00319822557503535,0.0056089264330812,0.00442063720789743,0.000920147590745213,0,0.000239528732159267,0.00387502412509044,-0.00217317058423616
"1496",0.00680818558479879,0.00887254434861284,-0.00106951586670578,0.00511284523721911,-0.00760156582070215,-0.00193121651470862,0.001242536417287,0.00310979879466089,-0.000904758729105781,-0.00181478263702284
"1497",0.00048787778525794,0.00439741898834844,0.00428258319773112,0.00300563191781222,-0.011610195307205,-0.0042378570972238,-0.00062050764099697,-0.000715019896269209,0.000724479350117102,0.00472724539946046
"1498",-0.00613200363417699,-0.00283304668914119,-0.00426432088874329,-0.0043799829704908,0.000734334038442697,-0.00194285646515402,-0.00667484386682349,-0.00548936684256296,-0.0084454905363941,-0.00904819863907314
"1499",-0.0037155668252471,0.00490696841170157,0.00535333509023461,0.00439925161765897,0.00749920570734997,0.00222467456402042,-0.00125025623533281,0.00551966631581902,-0.00146005966599916,0.0062089023060381
"1500",0.011752264763911,0.00429231761119886,0.00958454836427158,0.00253579684145366,-0.0149674489677191,-0.00527187923622263,0.00625868616620529,0.00811427190854497,0.00188872838942511,-0.000725868225068038
"1501",0.0111287508233366,0.00875389540443994,0.0150336004289042,0.00698597540359658,-0.0101848897272994,-0.00390604039610298,0.0102628733939376,0.00639225808861954,-0.0143517390616426,0.00254264592044251
"1502",-0.00742965383874417,0.000765692219063974,0.0157564548557665,-0.00045936475382502,0.00331894348700668,0.00140022712678878,-0.00140251929394708,-0.00352887400677682,-0.00240621912134487,0.00362325082674775
"1503",0.0057524854763138,0.00586557266224341,0.0134435247695819,0.00597575671077544,0.000165456092837912,0.000652814669569013,0.0113905819533606,0.0144006346534318,-0.0121219987368173,-0.00469318791637974
"1504",-0.00907704569098922,-0.00938099141641757,-0.00612251366755256,-0.0114233768959863,0.0109152267302708,0.00270171425250698,-0.00308542892556896,-0.00667216221186828,0.00375637647921812,-0.00181354069069395
"1505",-0.00308122912415942,-0.00204770051405267,0,-0.00208013281537944,-0.00179950045085542,-0.00102235866234912,0.00139233247805959,-0.000486944254985633,0.00180872573057145,-0.00327037887043391
"1506",-0.00421470108302857,0.00102591923083284,-0.00102679602599887,0.00301064514486016,0.00359689375220618,0.00205862387971223,-0.00494494053733108,-0.00097421959741284,0.000996164892173024,0.0102077748250822
"1507",-0.00134045107377812,0.00435560856149486,0.00102785141975192,0.00563561244552724,0.00335567415791393,0.00204448399545165,0.0012424920019718,0.00316869135752151,0.0023635091576284,0
"1508",-0.0108085609677842,-0.0142857351145594,-0.00718668069125394,0.00367456059826443,0.00570927820761602,0.00231892719849314,-0.00604940798692333,-0.00753133217874769,-0.00384717662330147,-0.00288700503424477
"1509",0.0169963533364959,0.017080901525145,0.00827296060123106,0.0148743293150688,-0.0172739087310653,-0.00527449165732941,0.00920743135202273,0.0122401185189969,0.00921895517959803,0.00542888193349578
"1510",0.0256303547444177,0.0145038868304797,0.0246152408856555,0.0196168539918598,-0.013368375253502,-0.00455826440702101,0.0162361099656938,0.0133007474614868,0.00709785194178858,0.00359966281133017
"1511",-0.00225922437972725,-0.0135441842167113,-0.00900886654513822,-0.00707668591585353,-0.0135493578666149,-0.00514041164752288,0,-0.0152746267665644,-0.0120733040641454,-0.00824960277536924
"1512",0.00439123332008196,0.0071193523126285,-0.00404032384835362,0.00200457270809595,0.00390006045792202,0.000469790829401795,0.00608643316778279,-0.00169642692131189,-0.00471460926888234,-0.00433994176907604
"1513",-0.00273240634739347,-0.000757474001746972,-0.00912786991947345,-0.00755715184280126,0.000422388868023482,0.000562835604980272,0.00151253363898785,0.00315602420433403,-0.00629524424962291,0.00181617565745906
"1514",-0.00287730503905614,-0.00202115842246875,-0.0133060400096615,-0.00895863156006316,0.00658467412160224,0.00244009026843317,-0.00196323994906156,-0.0084705299589064,0.00708778178269132,0.00253807371799342
"1515",0.00254189395144722,0.00101254725023914,0.0134854783237872,0.00429377552934795,-0.000922336827764103,0.000561733744737225,0.00378256835620161,0.00488155036257365,-0.000435930498703718,-0.00144667207169502
"1516",0.00794967642728239,0.0174508620240785,0.00818831246555196,0.00877579502143822,-0.00277066573603113,-0.00290052290240239,0.00241182048948541,0.00777264581036441,0.00928401117564914,0.00362186399421871
"1517",-0.0000678234501764186,0.00422568666636214,0.00304558934532562,-0.00803023368953037,0.00892349865889663,0.00319024226435061,-0.000150301249213003,-0.00385590536606195,-0.00567970133793549,-0.004330618978589
"1518",-0.000680322946384648,-0.000742631237166669,0.00607302399280218,0.00427242774722369,-0.00275332421427432,-0.000373705726234075,0.00150419667038082,0.00435494747022047,0.00298022479796622,0.00652420086718264
"1519",0.000680786100790698,-0.00346784947289625,-0.00301823885992192,-0.00425425176394378,0.00460212902649348,0.0024325896709092,0.00465529251561603,-0.0019273248145012,0.00631425680450537,-0.00432122496650611
"1520",-0.000136075672291569,-0.00472261916597283,-0.0121089677932892,-0.000899441775025323,0.00208149777319111,0.00130681506439245,-0.00104651230849861,-0.000482663929676108,0.000553617132795337,0.00108497613651792
"1521",0.00646004424102364,0.0107389030213154,0.00408572109101901,0.00562683649188767,-0.00997312808768624,-0.00456777565185951,0.00224449829188833,-0.00217346311735467,0.00430379358021993,0.00433527532181133
"1522",0.00223020868562207,-0.00222367201075802,0.00406943783372737,0.00223790411444647,0.00772324246046563,0.00280904975707208,0.00597177947661232,0.000967933329632853,-0.00159173547872404,0.00647484275670118
"1523",0.00539291292846622,0.000247174014537332,-0.0101318081786134,-0.00156315310792732,0.00191587118361114,0.000840797740921717,0.00504643717426156,-0.00338475763189894,0.00355633094748486,0.00285914600816461
"1524",0.00160940017237254,0.00049533330929763,-0.00818839847392483,-0.00536778776164171,-0.00149654763449525,0.000466397648563266,0.000147515067911552,-0.00388169743873401,-0.00281047843600513,0.00106912297437733
"1525",0.000267960849967386,0.00569163730380118,0.0113519086776011,-0.00359803148627846,-0.00349700967269806,-0.00167850523659485,0.00118112235354007,0.00487092210583073,-0.0109675199021344,-0.000711914167553562
"1526",0.00562235080346718,0.0135335892210426,0.00714302312084869,-0.00338527204206618,-0.0137047172010613,-0.00663339951364161,0.00412926664444413,0.00581665217061511,-0.00477018962669051,-0.00213755737961818
"1527",-0.00119859046771442,-0.00194200628675523,-0.0151974852360464,-0.00701984792885413,-0.00364288706347526,-0.00206853798819262,0.0010280861005052,-0.00578301438742579,-0.00224090266694921,-0.000357010471621177
"1528",0.00393153951192549,0.0051080634533851,0.0133742825737344,0.0111744319597393,-0.00552739717124573,-0.00150825884262806,0.00190728342384761,0.00290855799358947,0.0043671597140813,0.00571428109331551
"1529",-0.0039161430408261,-0.00121004045205442,0.0101521256252073,-0.00473599382619538,-0.00170995331505941,0.0005661829189747,-0.00922534561492727,0.00338290742559799,0.00745386025672823,0.0113635906775538
"1530",-0.00246515657979085,-0.00411920011734201,0.0020101936931185,0.00203925590258458,0.00488174200992497,0.000849447654696744,-0.005764330165558,0.00120478907646571,-0.00610398290765168,-0.000351118811761197
"1531",0.0102873016939256,0.0104623951558169,-0.00300896043819077,0.00655805944783805,-0.0129846381392362,-0.00339774865139741,0.00668972859530848,0.00384862479504333,0.00155086851521458,0.00386373583612265
"1532",-0.0112407869968901,-0.0276907951411364,0.00100582600776833,-0.0132554799283364,0.0128094014702196,0.00577649604456365,-0.00206734742995374,-0.013419725600041,0.00340664608374075,-0.00349897458315218
"1533",0.010098126330627,0.00693382650390384,-0.00301509348394391,0.00113862275635035,-0.00888744853401358,-0.00357779436811323,-0.00133203585313035,0.00607268905390601,-0.000246870370370411,0.00386237920578703
"1534",0.000728021823759306,-0.00270520300313681,0.0131049552968387,-0.00113732776907105,0.00819136020167033,0.00302398624199585,0.00177818070864699,0.00048253158881284,0.00265492702775694,-0.00139907150236718
"1535",-0.00132288322874541,-0.0120839783100902,0.00298498078161336,-0.00887961919340952,-0.00222354850189899,0.000470670847958488,-0.00473297301194098,-0.00627386383840201,-0.0033869265557418,-0.00385290912519543
"1536",0.00556415116120723,0.00848745669210804,-0.00396817589787246,0.00735124116409835,0.00385701363290147,0.000753566436811681,0.00995682751843918,0.0106844638707497,-0.00166824645744557,0.0038678114512305
"1537",-0.000197665293095506,-0.00594083461515915,0.0109562587997001,-0.000455972314978403,-0.000768314725543062,-0.00103458932168687,0.00102989653104379,-0.00336333040697068,-0.0115739921952223,-0.00350257911454177
"1538",0.00164742392437867,0.00821729990963527,-0.00689671159130822,0.00273777936484443,-0.00247816747835983,-0.00103633454010821,0.00587984308451439,0.00168725156398075,0.00118974329097821,0.00175744514794096
"1539",0.000854960143178651,0.00493953307451722,-0.00396817589787246,0.00500559372390064,-0.00813795832713815,-0.00348857384130374,-0.000438283393984218,0.00553566777858783,-0.00525358687381061,0.000350872390607826
"1540",0.000920206443347338,-0.00737317110848434,-0.00996003237449927,-0.00045266893267315,0.00906823442217664,0.00425741043092942,-0.00394758032801623,-0.00526567120131172,-0.00440111277457822,-0.00140306948977265
"1541",-0.00118218338712961,-0.00321840525930639,-0.00301823885992192,-0.00362389690537634,-0.00290982756995539,-0.000942321934421342,0.00117449973342687,-0.00433105995338157,-0.0163562418810391,-0.00421490567380778
"1542",0.00749483418278207,0.0111776513510475,0.0151362592043864,0.00204563882273856,-0.00497864472402565,-0.00160305134963878,0.00689029113190553,0.0113581206640634,-0.00276061256935711,-0.00388012635360513
"1543",-0.012463107901642,-0.0132650209435572,0.00298201355870753,-0.00884736093238669,0.00301951477936968,0.0021724799761893,-0.00844513458137131,-0.00740754576320146,-0.025043455545697,-0.0113313996413342
"1544",-0.00607924084443123,-0.0164301081760937,-0.0118928402111043,-0.013733219138988,0.00584834030764259,0.00197960915148099,-0.00778258883056493,-0.00698098047563001,0.00779181843909371,-0.0114613456196369
"1545",0.00977271623248188,0.0151863493206579,0.0160481635949388,0.00440936580270823,0.000684243054825728,0.00122274885219764,0.00858416169020648,0.0050904061790189,0.00229331680950451,0
"1546",-0.019026971124757,-0.0309151555772628,-0.0138204624801093,-0.0134010146933891,0.0196530710450555,0.00770387879659351,-0.0168748776354299,-0.0159187325090309,0.00895597170062135,-0.00471015522293972
"1547",0.00684544403100151,0.00694634947934181,0.0190193101774498,0.00562071025481359,-0.00578202183065024,-0.00186473829502742,0.00880599320731679,0.0137254369243522,0.0121809320249042,-0.00182014263204167
"1548",0.0125984658706324,0.0166070565570358,-0.000982553146880338,0.0109451962304183,-0.00295052119039829,-0.00046699354598434,0.00769337421006866,0.010880384005681,-0.0105619894343746,-0.00619988201925725
"1549",-0.00197510661325917,-0.00276472588357546,0.00393327931458254,-0.00460737606475814,0.00185998396148124,0.00140163519254166,0.000146962753838409,-0.000717626807934857,-0.0101572551523531,-0.00440368522061918
"1550",0.0032979724370974,-0.00453610714988695,0.00979419300730111,0.00231466402842639,0.00544565889099258,0.00249460648539546,0.00190832547445274,0.00694108961636952,-0.00366011764705887,-0.0070032599178137
"1551",0.00532529122050107,0.00405028336696289,0.00581962699019178,-0.00946682774455287,-0.00529842248940504,-0.00232985147575415,0.00747258775011317,0.00499150307261731,-0.000918387550270405,-0.00371197812652269
"1552",0.00895912301859791,0.0115987933786199,0.00192866963742588,0.0121210991744982,-0.00287479951450831,-0.00102765264655924,0.00770811625283896,0.00402068631077457,0.000525292176126957,0.00931452061308158
"1553",0.00136122108783265,0,0.0125121398270844,0.0048366404835305,-0.0090727497979588,-0.00317905875887037,-0.00375256815838576,0.00235574846562692,0.00557810061759745,-0.00553713659489818
"1554",0.00181229831602558,0.0067296159838941,-0.00950568692029896,0.00275032973802447,-0.00770226024555487,-0.00384641495001548,-0.00362160272962286,0.00164544590040894,-0.00352407501204921,0.0066815377053342
"1555",0.00426388714052295,-0.0007423231950483,0.00479840231925421,0.0086859105652628,-0.01043459411423,-0.00508511908209286,0.000581526344062056,-0.00351945766585926,0.000131017091741237,0.0029498120940703
"1556",0.00379548252274331,0.00322088848620661,0.00573039786134766,-0.00543865515573105,0.000958513024238661,0.000473330479054734,0.0039231998908793,-0.0014128106571677,0.00183352751728982,0.000735284073664522
"1557",-0.002243238381753,-0.00271656060786751,-0.0104460255871022,-0.0113922413851991,0.00722630302186689,0.00274348592981721,-0.00361832350716251,-0.00589492394392244,0.00784363004628963,0.00220426929571249
"1558",0.00141342130939615,-0.0024767863968812,0.00575789461573595,-0.00944896999905342,-0.00103714782019348,-0.000849394481487575,0.000290692915617452,-0.00047416694489355,-0.00343730457957969,-0.00513193244750831
"1559",0.00532391415555389,0.0139029491983944,0.00572543888202626,0.0041879403293934,-0.00302830765810913,0.000283767549480007,0.00537305624524298,0.0163741704167963,0.000130085900557519,0.00736920964057641
"1560",-0.00132041821934981,-0.00171404606597669,0.00948754324451229,-0.00903614187061463,0.00468657446721976,0.00349253371544078,0.000433352912377227,0.000280840070292943,0.00208229447277497,0.00219455661418477
"1561",-0.00551882051216079,-0.0139810268746577,-0.00469918787408674,-0.0112228861208624,0.00760217019462073,0.00329255510888182,-0.00274332209880179,-0.00726501873241892,0.0089610714285715,-0.00583944890513199
"1562",-0.00232322780448802,-0.0024877534779405,0.00566567584939914,-0.00709374777587979,0.00677293835548154,0.0030942943738812,-0.00709422501887358,-0.00613815343068014,0.00450506485696156,-0.0073420437609536
"1563",0.00698579332894567,0.00573588611663345,0.00751169327968682,0.00571530203891601,-0.0111557210614222,-0.00383267790611641,0.0058325319745447,0.00356324858527546,-0.00454899404729647,0.00702653066856218
"1564",-0.00854252931665189,-0.0116539504672987,0,-0.0101822082596474,0.00964504860719373,0.0026274596473943,-0.00333420194883161,-0.00591715257645398,0.00566393144313371,-0.0044069196129316
"1565",0.0080328056360095,0.0102863250640688,0.00372779200861206,0.00382805569890365,0.000767450608307074,0.000374866921649675,0.00610895132526368,0.0128571299408773,-0.00447998080000001,0.00184431274578434
"1566",-0.00417762882097994,-0.0156447353923791,-0.00928493298364697,-0.000953665609279675,-0.000937116753123801,0.000748072968238311,-0.000670473970156404,-0.00188037942732977,-0.00199291542283031,0.000736442796368086
"1567",0.0080030171277099,0.00479344453854669,0.00937195091986398,0.0143132823768057,0.00119401435426281,0.00102792569904842,0.00744070805188057,0.00894937150634223,-0.00334967781017526,0.00919792752690629
"1568",0,-0.010042983513997,0.00464246649182365,0.00376281881422691,0.00852114548665384,0.00429635713670073,0.00159326189819042,0.00396803843639804,0.00413650462683246,0.00510390617331535
"1569",0.00307317370959503,0.00710132900310834,-0.00184825011259038,0.00210875785732667,-0.00506950169080422,-0.00185987557195832,0.00462682684927507,0,-0.00585738925169044,-0.00943056091566707
"1570",-0.00395740249398568,-0.00528827752008343,-0.0388888045993555,-0.0107551799611744,0.00753147725490555,0.00265889618937032,0.00316642379940779,-0.0179021495649229,0.00142441569616869,0
"1571",0.00493470513786431,0.0108860310598162,0.0125237609887194,0.000472763324836922,-0.00405426792988539,-0.00195398162609495,0.00258260851995695,0.0187024499167037,-0.0144824790131568,-0.00476013385914431
"1572",-0.0101396775832862,-0.00500880786458358,-0.00380561130918033,-0.0118118593939163,0.0089899359169987,0.00419487497058113,-0.00529490313401815,-0.00720447416718939,-0.0111526410684805,-0.0169242426921778
"1573",0.00405872009532549,0,0.0410694342067128,-0.00286890444586307,0.0119356578008727,0.00399185928128221,0.0146739578076966,0.0203653572296267,-0.00291914689628192,-0.0011226621444842
"1574",-0.00449134621202563,-0.00604052030041446,0.00550464618904667,-0.00239767926295797,0.020184637936226,0.00314386262643174,0.00269389046133051,0.0142235006692617,0.01676761672349,-0.000749411160418934
"1575",0.00676770173031493,0.000759429565416969,0.0100364713533707,0.00168246587379439,-0.00765362721002194,-0.00322618773507055,0.00933271309790751,0.0022620012803205,-0.00425360911267092,0.00299958406858414
"1576",0.00345650219261318,0.00556682082357263,-0.00812985193100046,0.00983682720010215,-0.00246128244933197,0.000369735135919091,0.00042042084013616,-0.00112856390036864,0.00775494196227822,0.00635520752959895
"1577",0.0122488982984679,0.0158531062833767,0.0209469578512131,0.00950340336055233,-0.0137362171013132,-0.0041598445354577,0.00588151986209806,0.00610027591895923,-0.0168905443299999,-0.00222887210996559
"1578",0.00327716964248115,0.00569715269783755,0.0115968915374323,0.000941355151300449,0.00191827731824268,0.00111433511793724,0.00487246467816749,0.00381744297698261,0.00199006965174142,-0.00409532978060922
"1579",-0.00245006710222984,-0.000985175061679056,0.00176357180756126,-0.0152832982924004,0.0148993496764074,0.00556317967008835,0.00581892393587546,0.0123046167552618,-0.0470043419992517,-0.0123363959983461
"1580",-0.0231737033524951,-0.021943017563224,-0.00792250877471989,-0.0243554284379582,0.00869331285308439,0.0022128971020039,-0.024931462982469,-0.0227625116244619,-0.087808261642409,-0.0299015704037351
"1581",0.0147627866202569,0.0143688340997836,0.00976052563283747,0.0205582791888563,-0.00821171543102639,-0.00285174157235635,0.0158218767839973,0.0174127789445471,0.0113472319145111,0.0105344659073492
"1582",-0.0146112786542953,-0.0280818155904055,-0.00702993468240753,-0.0158273209691766,0.00664030850568609,0.00184516522327738,-0.0120987724459122,-0.0111135013193092,0.000527048180864798,-0.0146718133830123
"1583",-0.00625391736687242,-0.000766713416890719,-0.0070795310292503,0,0.00244333653013151,0.000552280991292564,0,0.000449210375425002,0.0107624599519254,0.0105799947329301
"1584",0.00869349579663004,0.00690879941571376,0.0106950995901169,0.0146199606928448,-0.00211260739108798,-0.000551976145359734,0.011543013895696,0.0146036357877208,0.00871182407940818,-0.00232653110253789
"1585",0.00443817227149279,0.00482845485276773,-0.000881946455283389,0.00480276969686333,0.000732960763767165,0.000552280991292564,0.00139157778762877,-0.00221415799482649,0.0179374989448771,0.00310924862864859
"1586",0.0103087259751244,0.0171979341299593,0.00970863969599822,0.00478015056031289,-0.00349810487100088,-0.000643868007821013,0.0058366949745341,0.00199683559687358,-0.00739658480333205,-0.00619922233375714
"1587",0.000634244593010536,0.0079560480107348,0.00611902462185365,0.0059467268251816,0.00253083762883,0.000460306510481123,0.00317760883716689,0.00442998009871576,0.0108853736526382,0.0109162716021534
"1588",0.00405355597589341,0.00518034496362296,0.00521308418961342,0.00898555656382349,-0.004315973857413,-0.00110487573591245,-0.00123980617057617,0.00308700868005385,0.0235600933569451,0.0131122044342977
"1589",-0.00176654709296309,0.00294467560774536,-0.00259292760324847,-0.0100772931387115,0.00916001917791465,0.00359455811234444,-0.00455022579622322,-0.00395653404562146,-0.00508367559543632,-0.00570989639238018
"1590",0.00669890406202045,0.014925363605681,0.00606563392562709,0.010416666086783,-0.00364721210552366,-0.000367674629913717,0.00775719807400588,0.0134626855133348,0.00986444511065376,0.0133996281898012
"1591",0.0023853186323135,0.000482107231851048,0.00775198436589664,0.0142926401100179,0.000569494162733886,-0.000183344600924396,0.00975919129093916,0.0041376211709907,0.00330288819459823,-0.00755569810693069
"1592",-0.00876703911121823,-0.00578291814946619,-0.011110921717332,-0.0108570306194804,0.0102734189087452,0.00326540549427468,-0.00680614779441568,-0.00303660408589379,-0.011627113213501,-0.0178911993642445
"1593",0.00928719371730891,0.00484710893249529,0.00432136847119646,0.00794004427338613,-0.00129050660872398,0,0.00383732293585659,0.00478567542277286,0.00574018137807242,0.0127906433562244
"1594",0.0101403684599244,0.0125421837559758,0.0137693800944205,0.00834097650208121,-0.023576983940432,-0.00852789645017138,0.000819398185035736,0.00974281663439869,0.00119784387257416,0.0110984797220384
"1595",0.00254071693292079,-0.00214395396871214,-0.00424449920910808,0.00137880293311099,-0.00248088837964111,-0.00129498192007804,0.00395645484623741,-0.00171536286996199,0.000422253513188808,0.00113548788016282
"1596",0.00506899315026166,0.00429697246314253,0.00170503193481375,0.00711327342421697,-0.00389601446910626,-0.00138868060164155,0.00584319748866458,-0.00536937753405287,-0.0124515587387221,-0.00340260002939397
"1597",0.00455068281307303,0.0125983699896208,0.00851052955441767,0.00774698344980873,0.00158107141862596,0.00120551730365759,0.00243188117125337,0.00539836338513355,0.0148169392072608,0.00455228966012333
"1598",-0.00281596878973833,-0.0103289045821874,-0.00759472229864255,-0.0072351616810703,-0.00257571543542112,-0.000185105764410887,-0.00512127796549045,-0.0124567820546512,-0.0115822611183781,-0.00037763835250948
"1599",0.00325392796454138,0.00403224380448708,0,-0.00774294546704057,-0.0107463955552783,-0.00565181298115636,0.00027075484493122,-0.00282781444177671,-0.00859308299968875,-0.00453344997004712
"1600",0.000795201072960161,-0.00496096164003212,0.0127549376839307,-0.00918099151653706,-0.00766313168012311,-0.00177029986104371,0.00148983585051199,-0.00937789806597511,-0.00838118158820145,-0.00455409573522136
"1601",0.0103341912567958,0.00189959912428939,0.00671717070042943,0.00463307243409328,-0.0108623876525918,-0.00401281505572082,0.0052739088557876,-0.00440335265544656,-0.00447876205556108,-0.00343117818564065
"1602",0.00538629211676556,0.00402806721669724,0.00917431085499154,0.000230509397574963,0.00669191261790258,0.0026236139907625,0.00887791703981167,-0.00309617408686491,-0.0230751980708975,-0.00229530155362823
"1603",-0.00469519320806189,-0.00330412694763427,-0.0148760734247843,-0.00345776562843436,0.0103970849555661,0.00476707979517643,-0.00319967752453409,-0.00155291133880264,-0.00401105979309735,-0.00115036996924256
"1604",0.0096769738490956,0.00710394124851632,0.0159397221604021,0.00439489566028972,-0.0126518073531896,-0.00539507819517382,0.00628653831321579,0.0135526159175514,-0.0225221052284915,0.0049904142640429
"1605",-0.000060177635464731,0.00352719315910033,0.00660572455265451,0.00253357763441753,-0.0011959449661314,-0.000748871736752532,-0.000531377980863668,0.00548007766011782,0.0308994261364461,0.00649353610594772
"1606",0.0014381008170139,0.00234276052210247,0.00574263848181289,-0.00206766149653614,0.00786876690834282,0.002621003667858,0.00465446680323467,-0.00893846216642336,-0.0165777833251103,-0.00569256107987448
"1607",-0.00741747208329024,-0.00864881063351763,-0.0106036819523699,-0.0110497629345979,-0.0148507972488316,-0.00793545020947539,-0.0247551741312482,-0.0217772157062301,-0.00707407408661687,-0.00458016862487476
"1608",-0.00289321267757925,-0.00495148563612136,-0.0420444234547276,-0.00744864294695058,0.0047378393290245,0.00103548929997821,-0.0139810413670317,-0.0179897836236305,0.0202364632372829,0.00460124309412979
"1609",-0.000845793722942023,-0.000710954894244442,-0.0180722511113149,-0.00867745451701907,0.00137189401597348,0.000376131435728455,-0.00385457173283388,-0.0137392650922583,-0.00631458282211894,-0.00381682028174757
"1610",0.00598861067331558,0.00497954730922046,-0.00613501345256218,0.00544146492904063,-0.0253426455805164,-0.0117462183508033,-0.00995042630236909,0.00371458225527932,-0.00201846598454203,0.00919547400448573
"1611",-0.0064944133211825,-0.00542694855753634,-0.016754710229114,-0.0127058556651978,0.0112440603288266,0.00408857055927569,-0.0199606329374151,-0.0168860293072748,0.0100381822594133,-0.00645409096761351
"1612",0.00369213621835596,0.00711742398013948,-0.00538129740529658,0,-0.00243204041274214,0.000094909751655825,-0.00954289702463451,-0.0115297565998537,0.013869279628135,0
"1613",-0.0143520074748168,-0.0209657834354084,-0.0225427453371393,-0.0181124453992463,-0.00339650295549243,-0.00274593998670636,-0.0122232406195177,-0.0211854185067967,-0.0203364964228931,-0.0118455806241523
"1614",0.00550630565567145,0.00986520465526741,-0.0119927239994686,0.0148057476525019,0.00529887647875071,0.00144515365032194,0.00247513317658155,0.00437747552266643,0.0193398823079434,0.0123741931688792
"1615",-0.0048068838890174,-0.00381218423484841,0.0289448557192795,-0.0121983256502034,-0.00923493407658116,-0.0025635426927525,-0.0116181288759271,0.00750615534345589,-0.0093765954646764,0.0038197756843481
"1616",-0.0140011107836227,-0.0150679839649517,-0.0381124450035611,-0.0179176600907734,0.0138058660214047,0.00485460875913701,-0.0107255972907712,-0.0206682136922014,0.00214455378672063,-0.00456618679793841
"1617",0.00905337852468624,0.00801330684387414,-0.000943304887089935,0.00838290043914336,-0.000607089561254992,0.00123131706043544,0.0187138468043972,0.00490816409944661,0.0074527373833313,0.00382265631848155
"1618",0.0127203319180036,0.00939523987563406,0.0387156940916444,-0.00513455630038273,-0.0178790177547936,-0.00775797602847783,-0.000583548178243021,0.0144074614222613,-0.0238042922713271,0.00228477333300514
"1619",0,-0.00167041700702819,0.0127272624954984,-0.0135168258615439,-0.00477210516642823,-0.00247868310206278,-0.00875247760626385,-0.0122769409982993,0.00495200333847534,-0.00379945755776012
"1620",-0.0103155939699208,-0.00980179458525787,-0.0197487024791646,-0.0189334553775744,0.0118983812782134,0.00248484223853063,-0.0153053561696114,-0.0216916755394456,-0.00515157525531462,-0.00877181068797406
"1621",-0.00827728666935157,-0.00120687914815021,0.00274747422721555,-0.00685637598720379,-0.0143032610865873,-0.00448093714677955,-0.0146464918474155,-0.00747345314050207,0.00750469043151969,0.00115427429577508
"1622",0.0152088105758315,0.0120858374007189,0.0237439842967693,0.0212219749922562,0.0156684130400886,0.00756656905048048,0.0304870108656301,0.0256020774277721,-0.00379884543761644,0.00653342551185299
"1623",-0.00627268546573745,-0.00740375542300398,-0.0312220024283051,-0.0157735313764443,-0.00236660767530794,0.00133021114446508,0.0025018747545773,0.00244731375173735,0.00515917432484025,0.00420005822399827
"1624",0.0077218656560798,0.00986520465526741,0.0267036217215912,0.00915752717963714,-0.00527136837631981,-0.00237317024450978,0.00132127551948247,0.00366206223651622,-0.00490953681742734,0.00228141593051934
"1625",0.00790545124827702,0.0033357648199801,0.0170402140782369,0.00428572360040613,0.000529897418121372,-0.000570806079848829,0.00161333177607648,0.00997306468299319,-0.0122598411524305,0.00189678735838483
"1626",-0.0138166327888394,-0.0189979924016292,-0.0123456942594019,-0.0308735922872415,-0.0103283963207428,-0.0137104376609838,-0.0300102438842902,-0.0236025300491807,-0.0116552557460359,0.00151455709395831
"1627",-0.0247783648131823,-0.0326796632709999,-0.0410715799651026,-0.0448070783973519,-0.0164122772845122,-0.00453724680902956,-0.0390887882309192,-0.0434139388238095,-0.0535262900230122,-0.0325141227318189
"1628",0.00321012503389451,-0.0090091098519387,0.0363129655027337,0.0143710768966903,-0.0169589663937518,-0.0105704709248188,0.0117795952027309,0.00489204857795089,0.0117314322286639,-0.00625247726745759
"1629",-0.0126357201452248,-0.0154040636190412,-0.0278526991760913,-0.0203152521688927,0.00415148933332588,-0.00244991237873871,-0.00636453298025585,-0.0190053490590819,-0.00895644120856198,-0.00432562145749138
"1630",0.00961397156877597,0.011864226597305,0.0129390192661356,0.0212823257454202,-0.0089112287364006,-0.00117873865017748,0.0184348217224202,0.0177812040804006,-0.00371176470588241,0.000789878627295737
"1631",0.00990133221143519,0.00726335777673537,-0.0045618070703537,0.0157625083989912,0.0064885246297961,0.00403245046220291,0.0149572800994002,0.010430091339747,-0.0420345181660766,-0.00276239324015415
"1632",0.00586947893275092,0.00463531628637681,0.0245786334757834,0.0200656334403804,0.0102228444690284,0.00538906908429526,0.0178489377690627,0.0198712071210956,-0.0197835392271182,-0.000395720742039196
"1633",-0.00409716764178403,-0.00666476159840501,0.00808644680784032,0.00574719525660794,0.00683771398616972,-0.00116969370323905,-0.00434671127718445,0.00961555232948785,0.0273417193834444,-0.00514652842086805
"1634",0.00585988950797867,0.011870818559782,0.012477470367521,0.00311710930183406,0.00201462908074124,0.00038113090806946,-0.00526838175600453,-0.00451131991465659,0.0169590796997812,0.00636692819458662
"1635",-0.000929835608377227,-0.0104564664297169,0.00704231870104732,-0.0178666387734877,-0.00063396238469593,0.000390377417186727,0.0116522207801539,0.00881172522619345,-0.00891599130477971,0.00395407799903147
"1636",0.000433705367698822,0.00128878180956504,0.000874079055664945,-0.00922745232310618,-0.00299106586794318,-0.00195241221124531,-0.00433810318969807,-0.00349394605683417,0.00574756337157267,0.00905876382185755
"1637",0.0107892837519714,0.00180184093462366,0.0131006125023372,-0.00638634480221745,-0.0340874635972368,-0.0168230870866967,-0.010516595573388,0.00776346752412627,-0.0219480043390426,-0.00234196863799574
"1638",0.00570459188211281,0.0107911329533872,-0.0068964459367834,0.00133884065020928,0.00969338937824182,0.0058698251431879,0.00394743529259611,-0.00422447443570417,0.0120247781192235,0.00508608309389769
"1639",0.00719712493363023,0.00279619751455162,0.00520800473925953,0.0131050755871651,0.00102510414207879,0.00168141064406901,0.0127045428339589,0.00798598209222812,0.00928793390866134,0.0062280993616175
"1640",0.00036331173984383,0.00709753154826909,-0.00345416716761626,-0.00950355991359875,-0.00782133746985669,-0.00355475000522598,0,-0.00594209620844754,0.00273581488801655,0.00309481492883301
"1641",0.0136209662566174,0.0279388308908901,0.0294629253595371,0.0490404529014179,0.0117306127861088,0.0100080983247939,0.0276283914297046,0.0328767427994021,0.0272013318032576,0.00501346891729848
"1642",0.000417981545569823,-0.00759079167776355,-0.00168343473365629,-0.0106707550785743,-0.000834838920382164,-0.000784962069088069,-0.00653964646933591,-0.00795752326318011,-0.000885391192617324,0.00383732509349644
"1643",0.0038208968143858,0.00444137163287217,0.00927472745469027,0.0102722151161614,0.00529159373827781,0.00314203351466391,0.00365662040868142,0.00607677540435358,0.000402827690393126,-0.00267588302880972
"1644",-0.003746813293524,0.00122804711819269,-0.00835419018936356,0.00406713733856279,0.00341670937027883,0.000489008483383513,-0.00160307479594168,-0.0026578324566997,0.00571749879207606,0.00114992905154732
"1645",0.0025668890230095,0.001472123069298,0.00926700892380716,0.00911408664055435,0.00184065331119676,0.00440249118018188,0.00525552022070319,-0.00314906988418795,-0.0125710546286417,-0.000765765091293669
"1646",0.00547763937209766,0.00857420628632366,0.00500828824877519,-0.0117913015954239,-0.0124930084062882,-0.00467552549714656,0.00624480235731117,0.00267326363411158,0.00559521569899446,0.00421458075059888
"1647",0.00177655214989292,0.00291486607056513,-0.00747509967911431,-0.00279245800647998,0.0158133184435079,0.0054805325079097,-0.00101061754369891,0.000969198458304676,0.00887024419207738,0.000763017835870849
"1648",0.00195082151427406,0.00484383371658526,0.00251053589092409,0.00992848278034852,0.00146536451002532,-0.0000972897861230004,0.00288930721992253,0.00508479973127218,0.0298137236846479,-0.000762436083540319
"1649",-0.00212368953689501,0.00168707286960923,-0.000834703068147924,0.0108394152000115,-0.00420612314908531,-0.00116801499004271,-0.000431916444538216,0.000481785201643214,0.00675264690321775,0.00152611420787818
"1650",-0.00366580019943052,0.00288742501182582,-0.00835419018936356,-0.0102243204883347,-0.012671723049273,-0.00672393427031914,-0.0194553870156247,-0.00866858387867486,-0.0171922278903276,-0.00799996926074609
"1651",0.00243284562661095,0.00575819445671866,-0.0185340178476145,0.00579476787041,-0.000372254333199207,0.00147124441329383,-0.00117582753394996,0.00364352898287068,0.0093347581737977,-0.00115205797759044
"1652",0.00106553351574301,-0.00238557661455485,-0.0231760362093831,-0.00225436029572368,0.00614020913104318,0.000882062925002591,0.00264886070286652,-0.000968036199426758,0.000854907917228864,-0.00615151468866593
"1653",-0.00307490346169903,-0.00382606153074738,-0.0219685093459978,-0.0125533149136662,-0.00730506038891876,-0.00205565986173339,-0.00792491857295852,-0.00823647325457566,-0.00240719057623229,-0.000386841912370151
"1654",0,-0.00336049437157837,0.00898469588742135,-0.00228829616458914,-0.000372509190053605,-0.000294018467300594,-0.00118361570941572,-0.00610635735291465,-0.00272441813089119,-0.0034830042132139
"1655",0.000712244199457146,0.00602120863363198,-0.000890250450023777,-0.00586142819093938,0.00363427537284222,0.000686968322919812,-0.0137736967453873,-0.00442366176214148,-0.00124879805060862,0.00699035586535879
"1656",0.0115577925816681,0.010054962329678,0.0276290661155072,0.0182002561563588,-0.0192680048092284,-0.00882602520218834,-0.00555647283147087,0.0118490250204111,-0.0105501563812922,0.00231393010372782
"1657",0.00169936229424339,0.00568870480925754,0.0156115795129477,-0.000251554209128702,0.011009536119658,0.008517870431485,-0.00437915882942874,0.00146340913089182,-0.00197456755410652,-0.00384769978730604
"1658",-0.00146224102504955,-0.00259264737108666,0.00256179911972887,-0.00629552256732846,-0.00769833863241565,-0.00314271835379432,-0.000606729115978588,0.000487289719014239,-0.00522320350408989,-0.00502117525665891
"1659",-0.00568282085975524,-0.00165410038256975,0.000851766862133063,-0.0126713438957371,0.00293322910305038,0.000295980203147916,-0.00349066197310954,-0.00146098121737848,-0.0137628961120818,-0.00815226196392715
"1660",-0.00324009855100482,0.00142049421957635,-0.0187233981143493,-0.0107802813121466,0.00745190942772056,0.00364371276482478,-0.00411227230007671,-0.00658355891554208,0.00145197223963889,-0.00665361032499945
"1661",0.00366462700526649,0.0103993119310941,-0.0052036824549595,0.0192010959459803,0.0027150365571289,0.00147203625934833,0.000917749127341771,0.0112910272634863,0.0218284249403395,0.0051221547324638
"1662",-0.00288553762906962,0.00163723509555469,0.000871719808036353,0.0020363936829253,0.00158754072728517,0.000686075874484215,0.00947283289575496,-0.00169863795738878,0,0.00705608126312685
"1663",-0.00118160296726522,-0.0037364830487272,-0.000870960574451574,0.00940071350650107,-0.00680600680197363,-0.00195855739232587,-0.00817305335441931,-0.00705125135301332,0.0178937725217267,0.0120669074580908
"1664",0.00295671792589847,0.00609457850795714,0.00871829225880649,0.0060406280622145,-0.0144560364663187,-0.00902681487376056,-0.0137341170966083,0.0017142128824168,-0.0107643998000311,-0.000384530976713426
"1665",-0.0051294363044897,0.000233194706378281,-0.00518569203136077,0.00325230491846584,0.00152421876418329,0.000891384507106796,-0.00216632644309733,-0.000978020277415448,0.00986380162617517,0.00807999927135161
"1666",-0.0139857377956232,-0.00512481718392477,-0.0139010809065686,-0.0114713589492452,-0.0135046038776172,-0.00553959589847053,-0.0189173922791649,-0.009052724211431,0.0208527286821705,0.0095419721382568
"1667",-0.0033057580568554,0.00210711028842137,0,-0.00857701291098423,-0.00347051574831458,-0.00388009753270291,-0.0230760984074047,-0.000740967597493425,0.00675829589553811,0.000378066669932675
"1668",-0.00639217591693753,-0.00887841594327454,-0.00264315294947437,-0.0188297739429646,-0.00870662682152457,-0.00429359587025258,-0.0135897958311434,-0.0113667498775476,-0.00429934372757068,-0.00113377136863213
"1669",0.0049158989064737,0.00353600211101202,-0.00883381801011862,-0.0018150859825169,0.0077097945604685,0.00541595078561197,0.0234541087628579,0.00324931768012826,0.00333309610382138,-0.00189184165773648
"1670",-0.00616010435930359,-0.011275508254302,-0.0142603531910611,-0.0233826276446367,-0.0109435741264207,-0.00628431540598096,-0.00208336707190926,-0.017438695237214,-0.00286893173731062,-0.0011372096858524
"1671",0.00911519019322271,0.0125921383894336,0.00632902662405876,0.0162274209284659,0.0101832844470124,-0.000401773701163899,0.00562075922432714,0.000506668509453023,0.00560302082818853,0.000379579586898826
"1672",0.00337230002905931,0.00610052696274477,0.0170710675216841,0.0117802395887014,0.0108559985927081,0.00562325329440361,0.0116575045587737,0.00734952830959124,0.0157367369284953,0.00796658499444414
"1673",-0.00372102854840117,-0.00629672190330932,-0.0114840496436156,-0.0108666256700494,0.00498561803710262,0.00199761520239594,-0.00378828342685544,-0.00654084946190403,0.00407711656384513,0.00564542635091381
"1674",-0.0160841623854406,-0.0194789642401143,-0.010723758423519,-0.023018751749978,0.012594486497606,0.00568083443951584,-0.00301083323521045,-0.015700085371021,0.00959765986558136,0.00973052179638567
"1675",0.00355114687253799,-0.00215424573837242,0.00271008288137375,0.00214199433965412,-0.00810350152972983,-0.00406307932783367,-0.004767824960069,0.000771668135262527,-0.000292453382084168,0.00148263579272623
"1676",0.00158601175114947,-0.00263834716267686,-0.00090122927633085,0.00801509299697378,0.00797994525036749,0.000994978704435212,0.00159674985412117,-0.00128518378685394,-0.00614448070359619,-0.0103626668671772
"1677",-0.003167646745316,-0.0108228040051618,-0.0198377868100197,0.00768583276967694,-0.00113108617935631,-0.00188883873255763,-0.00765275447270319,0.000514772241088313,-0.0091999708986521,-0.00299180861046588
"1678",0.00452187476646015,0.0143451350013324,0.0248391933574477,0.00631268217965886,-0.0141045777039981,-0.00567538138593704,-0.0083548058967835,0.0128635025918509,0.0133709929197368,0.00525124106240105
"1679",0.00827292725106199,0.00479390930415269,0.0152603063272101,0.0177729948509393,-0.00220674272996113,-0.00331019775829033,0.00712879814652423,0.00457172096021208,-0.0129012903225523,-0.00858201128343494
"1680",0.00126695274231259,0.000476704071525003,-0.00265257503338778,0.0118130846357691,-0.0139437180505793,-0.0076487253265185,-0.00852655757064125,-0.00176975985197381,-0.0182682825406718,-0.00225815504595728
"1681",0.00048213884927728,0.00643819916151056,0.00354620616787393,0.0147209536058661,0.0049734598438731,0.00608571703363792,0.0183355112233075,0.0032928637354348,0.0147503558566646,0.00565820345158907
"1682",0.00957624337669349,0.0106608078066182,0.025618281646179,0.026263097958052,0.000485505828788035,0.00201554895172573,0.0197576870076617,0.0217115544546453,-0.00178896765362513,-0.00637662282010609
"1683",0.00739691413382504,0.0128926632974826,0.00775195530259243,0.0075552527566416,-0.00698366248423921,-0.00462742090114954,-0.00124972569295245,0.0113662142541457,-0.0162049057962839,-0.00906001565387571
"1684",0.00313865535035784,0.00740543230994217,-0.00683757432136944,0.00072581937360594,0.00888874106535575,0.00505337991878063,0.0068835199853714,0.00464233047708573,-0.000303689073034463,0.00152390635694055
"1685",-0.0026564870137481,-0.0041350584581612,-0.00688474462277688,-0.0116026673814873,-0.00135550008496821,0.000100491159593874,-0.00637036450853989,-0.00583667761465434,-0.0305998412437321,0.004944778001164
"1686",0.00224889376965431,0.00392176664646882,0.00519946345052125,0.0066030715683254,0.00387789958094631,0.00130682844496932,0.00218897405224583,0.00660488317782115,0.00117491973329531,-0.00302796768043412
"1687",0.00578772244913717,0.0059743666387746,0.0129309172751784,0.0111759355918934,-0.00666378659833144,0.00220960358968769,0.0098299972529996,0.00801940460271089,-0.0107182209356907,-0.0125284973465647
"1688",0.00446250073667076,0.00137035206589675,-0.00425532854219601,-0.00216236285765947,0.00826369967212637,0.00200394783908608,-0.000772540223466733,0.00699151233705009,0.000395436940975102,-0.0103806785639978
"1689",0.0115742263485263,0.0253193403241885,0.0307694420025331,0.0418973759657824,0.0123420113790984,0.0124000855752158,0.0349465611672539,0.0277709823745171,0.0435572727272728,0.0217560449952168
"1690",-0.00167589229408016,-0.00489440656728224,-0.00497527314085811,-0.00531543800125811,-0.00590470705054269,-0.00345701638264095,-0.00388471875678087,0,-0.00196950996021172,-0.00380226857225308
"1691",-0.00699141655414948,-0.00558921221380415,-0.00833339782756015,-0.0223047260652635,0.00526952264034142,0.000991363854472072,-0.017248961675276,-0.0112543001163529,-0.0287666110056927,-0.0091603372497493
"1692",-0.0046277079315209,-0.00382172618226362,0.00336137545819759,0.00356455930007638,0.00733893991133749,0.00376267984435685,-0.0064103215990976,0.000236750347167414,-0.00320409505473651,-0.00731889206234926
"1693",-0.00235377148958393,0,0.000837476061017473,-0.00852451206671001,0.010785981772595,0.00364982815281567,-0.0066051048279403,-0.00189658378360791,0.000862414719033699,-0.000388042802127453
"1694",-0.00289026712918283,0.00225679380090948,-0.00251034918366,-0.00764284057249598,0.00205971477007028,0.00275212021271876,0.00343376256625572,-0.00237522603540463,0.00885155071748245,0.00155269384311052
"1695",0.00384541725770338,0.000675647599270857,0.0159395142673557,0.00409148021555161,-0.00700611126399087,-0.00215633013704097,0.0060664194636284,0.0050000521290976,-0.00776451630057939,0.00775195220958547
"1696",-0.00459677937455771,-0.000675191407817133,-0.00743170667447846,-0.0117449061907059,0.0024460241931632,0.00137506926908348,-0.00371057239709538,0.000236866172109274,0.00923389929388918,-0.00499997149863052
"1697",-0.00532815072693815,-0.00653009372406355,-0.00831955414839169,-0.0113996088538942,-0.00150154352088194,0.00166770962753926,-0.0100869952976603,-0.00213173278192802,-0.00612551751472812,-0.00425197135461264
"1698",0.00791628691890933,0.0077060385845118,-0.00419461640629648,0.019872391632223,-0.00303463311660324,-0.00222633565531993,0.0152062365655026,0.00688366265922769,-0.0280074675928559,-0.00659936835062425
"1699",-0.000944789851389904,-0.00134917510890986,-0.0050545356307804,0.00384884583478473,0.00151250250800028,0.00167111600569303,0.000617584978226837,-0.00117870460813696,0.0198250427747024,0.00976938764059976
"1700",-0.00922117710203973,-0.0049549256774819,-0.00762086377472204,-0.00383408901724047,-0.00160445759027705,0.00137372220108922,-0.0154322680327922,-0.00873274804405089,0.000944451455130668,-0.00154804612847681
"1701",0.00757696023545895,0,0.00170639302951736,0.0129899209935695,-0.000756238359669537,-0.00274366417018179,-0.00360479119416279,0.00309520362736482,-0.00511087435131308,0.00310081279751295
"1702",-0.00864507143029036,-0.00520603332571412,-0.0187391560374177,-0.00854877840244794,0.00406735000002922,0.000883698697368596,0.00440473247765705,-0.0113930750967044,0.00877262316266991,0.0069552021763386
"1703",-0.0116463483073648,-0.0102390749117928,-0.00347242279153903,-0.00958083802375642,0.000283257751080068,-0.000490190289120451,-0.0114332185760031,-0.00384177943755915,-0.00188026482200143,0.00345352149477884
"1704",0.000725063839531526,-0.00275854150382659,0.0235191423048662,0.00749678384313457,-0.00800632957951131,-0.00176858633058341,-0.000317040761872001,0.00964100462357553,-0.0101255963873533,-0.00726575415014186
"1705",0.0215577920097929,0.0205162825326919,0.0144681645147799,0.0235238998859493,0.00161437701676492,-0.00216492116818445,0.0239302781282804,0.0181426356770873,-0.0145904685227938,0.0127119685621264
"1706",0.00644297963363383,0.00609901695629111,0.00167778572994681,0.00445592707483389,-0.000284484576321464,0.00147940383782208,0.00959649283391628,0.00281367658351939,-0.0134384730048719,-0.00532534128258155
"1707",0.00399443174813885,0.00291862484155736,0.0016753258492892,0.00583713517160067,-0.00806015380538672,-0.0033479991667088,-0.000306884355197545,0.00327347949228995,0.00187605223288823,-0.000382403970200285
"1708",-0.00725434260808344,-0.00268618093017825,-0.00836128995790331,-0.00974932290532182,-0.000668711095783703,0.000197611323930591,-0.00322048166671773,-0.00838954737370112,0.00732720821741917,-0.00344303107689314
"1709",0.0139662733721264,0.00718298752000224,0.00927472745469027,0.00796985189982191,0.0125309454282911,0.00484013195055066,0.0181537366807185,0.00846052736886871,-0.00153561784040357,0.00767759687630321
"1710",0.00668319050226729,0.0147092350693416,0.0083540270934872,0.00627906007062462,0.00906961409686491,0.00570259236955861,0.0154126410519813,0.0139826347196401,0.0314068072575133,-0.00533326056285455
"1711",0.0067542596613257,0.00636913768189529,0.000828640986036078,0.000924441491199968,0.00215321459760776,0.0000967767269988151,-0.00193448424678799,0.00873360010287061,-0.00447339514163236,0.005744925346165
"1712",0.0000571243446967351,0.00152785657485222,0.00082788564691838,-0.00161599041134364,-0.00317662682154563,-0.000683975140771231,-0.00521850233438037,-0.00273424850036352,0.00102487191209888,-0.00228489091290041
"1713",0.00579178293304716,0.0126389559067939,0.00496281275683508,0.00971281725591333,0.0111528114745192,0.00694471559711141,0.0106416746598803,0.00525516453619557,0.0185855484662416,-0.00114502251469084
"1714",-0.00478904645371869,-0.00602552354044406,-0.0205762664843243,-0.0233621707941767,0.00389285505095915,0.00174833213670245,0.0020761873711399,-0.0065911371766455,-0.00502546791481284,-0.0152846645628761
"1715",0.00332233010547278,0.00736090370066944,0.0100842201204658,-0.00211077248661118,-0.00387775949532143,-0.00203630664343069,-0.000740030206492825,0.00205886833483948,0.00940237766100904,0.000388042802127453
"1716",0.00456774084470779,-0.000859679208255915,-0.0149750025661954,0.00470050302647995,0.00370792435523604,0.00174900831405989,0.00977489447745161,-0.000228267628651024,0.00431110874416207,0.00310321811263736
"1717",0.00159131936619339,-0.00408693751041977,0.00337831447686243,0.00584784098228863,-0.00341717455396395,-0.000969755866218724,-0.00689374008633714,-0.00411021443991255,0.000766449445307904,0.00386688312838346
"1718",0.00533384656839231,0.000647962351004061,0.00757567932269154,0.00325579393222819,0.00129722823609857,0.0013587079515831,-0.00841798368396673,0.00114627739346673,-0.00605081197994506,-0.00269645895743109
"1719",-0.00496718223225789,-0.00366933040288631,0,-0.00556325592263074,-0.00601530259255079,-0.00261740815370293,-0.00729813936475987,-0.00847423350418852,-0.0013099945654621,0.00308999375752017
"1720",-0.0028359459901649,-0.00498254130068621,-0.00501265856996591,-0.0102565326093236,0.00214178525415387,-0.00116651295730996,-0.00720183391016938,-0.00323415724267617,-0.0143519129158065,-0.00847131645656707
"1721",0.00238924637505122,-0.00631377618113982,-0.0109150816055275,0.000471270793460654,-0.0108243744619569,-0.0055464524710418,0.00634706807881646,-0.00324485058598456,-0.00618444506316651,-0.0124271349969011
"1722",0.00351834685037899,0.00591575149502455,0.00084896928915934,0.00612071137083592,0.000941240973721724,0.00196039016055294,0.00135168942943009,0.00279005913253672,-0.00110278852546963,-0.00432562145749138
"1723",-0.00316679435948186,-0.00936624848701895,-0.00848166358739999,-0.0201218851108377,-0.0119481914944916,-0.00449975665964475,-0.0151470387093249,-0.00765108198120901,-0.00197145338650662,-0.00276465649222335
"1724",0.00510577551639901,0.00945480453569636,0.0136866527032036,0.00310400648183951,0.000476377299988284,0.003045828867978,-0.000152040393290642,0,0.00505688219116451,0.000792149946476695
"1725",-0.0126433662595697,-0.0154650847580077,-0.0185653011413589,-0.0180906698654403,0.00847037365873948,0.00264547981655205,-0.0121843029453025,-0.0135515048996323,-0.0081760457903155,-0.00712309554301804
"1726",0.0134914646261726,0.00553098619782277,0.00773864754757136,-0.00218212373515103,-0.0240659028069679,-0.0112371137418207,-0.0134131015266067,0.00450051367792437,-0.0149017512713459,0.00557991813609582
"1727",0.000168971052433076,0.00308026807740225,-0.00170660719721494,-0.00510188287035085,-0.00377126216850021,-0.000494168207087919,-0.000781654041241642,-0.000235952203057388,-0.00329897009413405,0.00435987023310913
"1728",-0.00203035787086903,-0.00592242698366563,0.0128204935674774,-0.00537255398059033,0.00465924549640362,-0.000889784828760343,-0.00344074386804283,-0.00165076852735579,-0.0114636793865259,-0.00670879114630474
"1729",0.00802445720288403,0.00441321259197447,0.00759497722542379,0.00171889510451795,0.00367150940023064,0.00415645942234888,0.00706216315720321,0.0011810070621312,0.00326664769130214,0.00437042702655299
"1730",0.00498963158601162,0.00241657260942274,0.00837518105333612,0.0161762336318678,0.00616084375380765,0.00482883299364056,0.00794779549376567,0.00802249942240563,0.0115588036069809,0.0043511245202319
"1731",0.0043508439605775,0.00416367142536878,0.0141197022190696,0.0190546835457068,0.00200947598246648,-0.000784239862088976,0.00247363504136566,0.012406456879863,0.000402373873075623,-0.00157540193747197
"1732",-0.00349922485791498,0.00240083041547168,-0.00163818784902714,0.00899395166185646,0.00601557979640943,0.00353321926805794,-0.00694011598544542,-0.00346825356780556,-0.0114221203346203,-0.00670606351599057
"1733",-0.00217355282844089,-0.00239508023399848,-0.00574226492994034,-0.00609906649285885,-0.00759317337379972,-0.00371660629837167,-0.00760999234135629,-0.00719252347705712,0.000406794134958588,-0.00158862234773016
"1734",-0.00312778323306373,-0.0104757655763578,0,-0.0136886518421394,-0.0170235386543217,-0.00549789769550701,-0.00876358705128566,-0.0100492354256175,-0.0230174385445491,0.000795534102772777
"1735",0.00806830117212121,0.0099251746002309,0.00412551350889157,-0.000957291598718601,0.00165372225236227,0.00088873938149292,0.0053678115028355,-0.00165205656538103,-0.00149850978608446,0.012718632235597
"1736",0.00500266596514765,0.00502288076031876,-0.000821763131194642,0.00718552428310293,0.00932535689382985,0.00285973444387033,-0.00298360554639521,0.00118192037635145,-0.000166783388914737,0.00313971495238485
"1737",-0.000995434739305412,-0.00173867626602964,-0.00740151505925235,-0.0128418351666986,0.00288654770259389,0.000787419381292676,-0.00425263518226837,-0.00661307673897971,0.00450301041532697,-0.00117365263192004
"1738",0.000276828226068782,0.00152386593182774,-0.0041422113558568,0.00337277231747435,0.00374275464170437,0.00216137608924849,-0.00284730038558278,-0.00071316691543144,-0.00531295870258142,-0.000391771302957644
"1739",0.00243515255441307,0.00369506189916069,0.00415944063810203,0.00648238730173745,-0.00172024813274718,-0.00225499494452974,0.0103110098273143,0.00499634605324895,-0.00300451510599231,0
"1740",-0.000662649913939495,0.00346451567447392,-0.000828178858443662,0.010257652593576,0.000286551120870948,-0.000589693266329627,-0.00926383719888724,0.000473633823036002,0.0103800268741003,-0.000391844188296631
"1741",-0.00259654563300959,-0.0079841921630357,-0.00248772907255601,-0.0210152931538338,-0.00777805762304506,-0.00429452246832507,-0.00522968904510679,-0.0134881818142905,-0.0258491721420673,-0.00117599337105756
"1742",-0.0043205732254501,-0.0100066632034558,-0.00415626185096463,-0.00337653205537602,0.00367762868771848,0.00178068415817823,-0.0011152023266543,-0.00407763962492658,0.00323181658051008,0.00588701097795474
"1743",-0.000111429152028886,-0.00549331104861084,-0.00751256041295878,-0.00121021856871451,-0.00954599239559395,-0.00454209037258491,0.00223289478276567,-0.00192673157224277,0.0169549001098246,0.00195089246041613
"1744",-0.00439572385621689,-0.00397700098042242,-0.00841030673879595,-0.00581533427247749,-0.00282309438597272,-0.00248008102442865,0.00111379557727354,-0.00506748159894321,-0.0138379127529001,-0.00116836855358804
"1745",0.0111772521378701,0.0135313631078746,0.0127225308637888,0.022178854524078,0.00478373397505427,0.000895034482363721,0.00778916805380292,0.00654847818282422,0.00211327129044969,0.00350880445250534
"1746",0.0025422485029869,-0.00043766241451304,0,0.00143064980150509,0.00233163262774694,0.00119234228981036,0.00646674997355223,-0.000963985748440144,0.00986923635927694,-0.00349653579214948
"1747",-0.00358340289867043,-0.00394111175425071,0.0016753258492892,0.000476211199045062,0.00717365056579333,0.0041673023437796,0,-0.00241175304635033,0.0175409203346064,0.00311894620786823
"1748",-0.0112305714264259,-0.00681475179829194,-0.00919764514689414,-0.022132300224584,-0.0076995136593595,-0.00385409761744293,-0.0216266506538236,-0.015957641970949,-0.0078804711869972,0
"1749",-0.00330151366270537,-0.0108455808208957,0.00337555850871962,-0.005840921687015,-0.00378301085591437,-0.00287665428076778,-0.00672746830737503,-0.00491350586573314,-0.0212642725362876,-0.00932762588406888
"1750",-0.00011214624839595,-0.000447672980687708,-0.00841030673879595,0.00244805865204678,0.00486816064325901,0.00149243617401629,0.004031500703221,0.00197486599288199,0.0092146080884723,-0.00392313431467806
"1751",0.00623174669050774,0.0123126206365936,-0.00593724730411982,0.00659350911187762,-0.00368164080898581,-0.000496737375843326,0.00112425443240594,0.000246557438666972,0.00259679182267036,0.00315080387494393
"1752",-0.00318034728611272,-0.00457718604355328,0.000853196514758681,-0.00873400335598784,0.00447351182334366,0.00318039162241024,0.00529450143503563,-0.00813011005727615,-0.00868911339812661,-0.00471136123717364
"1753",0.017072743729412,0.0156251078852927,0.019584299178977,0.0199042794168083,-0.00503482338733252,-0.00376538979997854,0.0175551093164603,0.0116743143901157,-0.00876528430231294,0.00197235968110299
"1754",-0.00115591509022661,0.00307700773048181,-0.00842454067834442,-0.018401919110586,-0.000972311549765958,-0.00417660468025327,-0.0122334272639365,-0.000491192947463137,-0.0237224808798361,0.0023622536040393
"1755",0.00581692670129286,0.00328654280678453,0.00339849836177897,-0.0014799047874775,0.0153885706157386,0.00309605578192551,0.0077801810560818,0.00326201663633063,0.00975441560703727,0.00785547348507354
"1756",0.00534256615792605,0.0109194320079848,0.00931394075123526,0.00741103057075332,-0.00565966798217044,-0.00318630728393665,0.00141526457743879,0.00825438623348229,-0.0031913230431031,0
"1757",0.002191481268212,0.00691292488367923,-0.0134227910506861,0.0058854289698691,-0.00800660787212237,-0.00389511672936638,0.00174717572207039,-0.0017367025842262,0.00458594791035738,0.00311765026524369
"1758",0.00508389793794373,0.0049345193538457,0.0161565787917108,-0.00853263674044324,-0.00385363914485148,-0.000863483279778476,0.00110954761390047,0.00372793502720858,0.00551248932838044,0.00155406033549488
"1759",-0.0000545536473828268,0.00533745618857928,0.00502085729240598,0.0154904607981052,-0.00284082654219653,-0.000603629469462019,0.00126666058939806,0,0.00325513968228774,0.00271524598323292
"1760",-0.000162918778496057,0.00339754877048226,0.00915902312296324,0.00435834926303369,0.00687566907989168,0.00271595126579482,0.000790975103209357,0.00940803070394436,-0.0147712086380325,-0.00580270831542484
"1761",0.00473274033179849,0.0042329136681909,0.001650167202357,0.00771474783177206,-0.00634090477975613,-0.00451383486821177,-0.00316044925240555,0.0105468354667746,0.00632640615587476,-0.00155639897877735
"1762",-0.00958362792138823,-0.0229715852671426,-0.0164744407649028,-0.0385168944999583,0.00304326900437935,0.00392973904548732,-0.00158538684788301,-0.0189319443849404,0.0161901218690117,-0.0144193330254777
"1763",-0.00016393423906147,0.00086289235512349,0.00586263099452333,-0.00174158197225138,0,-0.000602196438151514,0.00587488009178716,0.0054427189813,0.0109322118644068,-0.00632664688813733
"1764",-0.00289802960681274,0.00172414058006032,-0.00333058529143804,-0.00947157438372137,0.00420883358259272,0.00281203083676407,0.00410419564264575,-0.00344440640572108,0.00176040739575489,0.00119377599891823
"1765",0.00614188064068544,0.00709978677970757,0.004177184416571,0.00427759820362161,0.00253401536527531,0.00160274746178191,0.0034584283492376,0.00172841592467576,-0.0056903765690377,-0.000794901731337117
"1766",0.000217714865813345,-0.00170914247444398,0.00166398773193044,-0.00325715299083518,-0.00272178728541139,-0.00490010903869154,-0.00156653842328036,-0.00419074961796062,-0.00589123884867859,-0.00954649111203931
"1767",0.000653966302452957,0.00085598260708708,-0.00332235499222389,-0.00527911547191251,0.00584892467121589,0.00261301161691518,-0.000470905740772576,0.00173276452052984,0.00287839477958696,-0.00803205995609246
"1768",0.00272290892950466,0.00962169761080922,0.00666676739170624,0.0176901508105338,0.0119207945705821,0.00841814288553722,0.0119309261724834,0.0071658313116485,0.015195027985776,0.00647764372042814
"1769",-0.0133050347694864,-0.00847107664299884,-0.00662261595163216,-0.0119195879479651,0.00498060279051793,0.00288241181127402,-0.00651551865263789,-0.00662411011825814,0.00631959909663071,-0.000402247119002164
"1770",0.0108975461883276,0.0128149281066674,-0.00250007237209426,0.0108069848753833,-0.00457478890845464,-0.00376595281165515,0.00624612467555985,0.00419868390632216,-0.00933728332516814,0
"1771",0.00539003183272557,0.00421784084912913,0.00751878395228411,-0.000248832379366237,-0.00105303553881309,-0.000894948141112906,0.00465550465173115,0.000245436390118314,-0.00191838353422624,0.00281690432515114
"1772",-0.0012994747320253,-0.000210046868007741,-0.00331666226867233,-0.00547121296449349,0.00670929967956813,0.00278809133128921,0.0023169656813582,-0.0012292651351844,0.00108638639189751,-0.00160515579427789
"1773",-0.00422973178103048,-0.00483107775260194,0.00249598159789577,-0.00500135988420125,0.00418814409139578,0.0023821187746198,-0.00323628916685315,0.00221580881069516,0.00951664571736677,0.00120581268813291
"1774",0.00294044036618102,0.00548745499420833,0.00165956913683796,-0.00150768384908495,0.000758722205690621,-0.00108948682895715,0.00695718696640824,0.00343903584791239,-0.0101711982138428,0.00240863827526017
"1775",0.000651808739510207,0.0012594481437902,0.00248564208992175,0.0133398843494583,-0.00246288107349824,-0.00277634068839672,0.00261042513126308,0.00416164771635552,-0.00426060996476041,0.00480578379051
"1776",-0.0081934249706026,-0.00167684792714884,-0.0198347796369822,-0.0245901379436451,0.0141497545556009,0.00676161506767081,-0.000459426969662502,-0.0107266606576381,0.0218139018069652,-0.00079720148395801
"1777",-0.0213359386010772,-0.0317095155849295,-0.015177037862705,-0.0262286155793848,0.00646169312686529,0.00404941906540524,-0.014708322432753,-0.019713935913466,0.00410542734128061,0.000398959814302602
"1778",-0.00491894635001366,-0.00542195751153829,-0.0128425523716129,-0.00392258965925674,-0.00697846567547211,-0.00304972908489476,-0.00606411623686165,-0.00351936432901567,-0.01087580332917,-0.00677829885603132
"1779",0.00595456836957142,0.0109029517490364,0.00867315816534742,0.0063008289458355,0.00243604828200361,0.00148019966244783,0.0101686302895325,0.00983867282343742,-0.0000826884927470628,0.00481735918529047
"1780",-0.00960502144994169,-0.0138050005585461,-0.00085989383194629,-0.0143489378831693,0.00822565301227374,0.00472915024452969,-0.00464605315305067,-0.0102426433947256,0.0125672099024525,-0.000799030209567286
"1781",0.0106003296935708,0.00393688207808829,0.00172098191777925,0.00926414936904707,-0.00287446485866805,-0.000980528900917599,0.0121364777301629,0.0070672969896397,-0.0220462478807361,-0.00399842815131779
"1782",-0.00585836720011201,-0.0137255403683397,-0.0266322684308478,0.00157353201458554,0.00669389712334567,0.00392614349174458,0.00307429630395051,-0.0105264103327246,0.00267177931047291,-0.00120436045501515
"1783",-0.0225053224114855,-0.0203223855833857,-0.0203000183109309,-0.0282797407535842,0.0121851853334913,0.00543607112597622,-0.0145592154493798,-0.0167173142460026,0.0102423519108119,0
"1784",0.00700478228474677,0.00901915347153315,0.000900951943294759,0.0202103493329646,-0.0106113132493998,-0.00301991178334038,0.0104200764882825,0.0118495333213144,-0.00272009561490272,0.00763659306640951
"1785",-0.00125457396350859,0.00402235310248633,0.00180018226054357,-0.00369785978516191,-0.0092454843722265,-0.00361533452977469,-0.000308168643813,-0.00152750368888532,0.00247956860037313,0.00199447064194791
"1786",0.0131873914004634,0.0213666596331767,0.011680133409929,0.0209435262923812,-0.0042927991390932,-0.00186296707299505,0.00739038630455036,0.0137684572353425,-0.00041225986963267,0.00398087837775551
"1787",0.0123953588661736,0.0124210527091853,0.0159857612847489,0.00571297542700222,0.000843418361313297,0.00265243034169393,0.00672484945912011,0.0125755490288733,0.00767073585732003,0.0114988169728101
"1788",0.00183683556117731,-0.0025830529991272,-0.00437058658356493,-0.0111025213555596,0.00280939585086015,0.000490147323370271,0.0091088531175747,-0.00571264288894069,0.00613898675843472,-0.00548796906493509
"1789",0.0109440148393729,0.0151059226274584,0.0140472573041486,0.0216709334918188,-0.00578942233733726,-0.00440719941171608,0.00346005670932481,0.0174868516757807,0.0117149611408225,0.00512409213369813
"1790",0.000494524872734825,0.00276355832755626,-0.00173150827647783,0.000255734473021629,-0.00516560569573732,-0.00236115226211142,0.000599986933029539,-0.00147367580602142,0.00056287390991594,0.00196075756439518
"1791",0.0051628133075885,0.00678408610314674,-0.00867296610869961,0.00102194176163151,0.00566435263617215,0.00473339155943342,0.00389541922355341,-0.000491408879728317,0.00851882986418051,0.00547949829681849
"1792",0.00551870380595343,0.00547443779004708,-0.00437460389881028,0.0122510750930569,0.000563541627052189,-0.000687512710751514,0.00402983426723003,0.00369005794983024,0.0132281777548517,0.00350334094595328
"1793",0.00119545308102165,0.00607363876747669,0.0219685905996063,-0.00932943348398396,0.00225179425382271,0.00245541531934745,0.00594636713591767,0.00955870563112704,0.00196618164425977,0.0143521342519306
"1794",-0.00662163812340089,-0.00666130202284876,-0.0120379662322032,-0.00687182440468903,-0.00421287029250439,-0.00195934977048529,-0.000295513561339611,-0.00242756035370528,-0.00886974083406999,0.00267682779140133
"1795",0.00590108908062636,0.005867646836893,-0.00609214160613236,0.00358792898912297,-0.00244396203869246,-0.00107974853788029,-0.00177404061706032,0.00803129860201968,0.0105329930434701,0.00190703312623652
"1796",-0.00114083518878072,0.00166677008669791,0.00788079885139448,0.00689463565862325,0.00527709315986402,0.00127776278099789,0.00162891235375429,-0.00193173865198537,-0.000156708466406141,-0.00266463921158044
"1797",0.00554684564113916,0.00665558424633628,0.0112944209221832,0,-0.00253088959225101,-0.00098156653693271,0.00162647144720474,0.00241912589262228,0.0110519123522197,0.00419845517025497
"1798",-0.000378768973002819,-0.000826447539567288,-0.00343624069655668,-0.0114125599908063,0.00892854204048654,0.00343807872017798,0.000442605220040138,-0.00241328784550887,0.00170557400939697,-0.00456098027062002
"1799",0.0000543570349351707,-0.00475615385528327,-0.00431051710861896,0.00076971312224261,0.00530968434880275,0.00293691636789828,0.00280311582355708,-0.00362850186583852,-0.00851331894131058,-0.00267273931650935
"1800",0.00524748393208418,0.00540214565955122,0,0.0189692072949168,0.00546740655253997,0.00117151680948657,-0.00102966669257598,0.00194221887750778,0.000702490042131743,-0.00306282394495516
"1801",0.00252921357167435,0.00289296453229371,0.00519483638109541,-0.0067924178049279,0.000552708157334658,-0.000975409038461716,0.00662718294596409,0.00508847148213265,-0.00452413427123555,0.00345609488391885
"1802",-0.00703195248814703,-0.0247269918199318,-0.0232556786659353,-0.0177303634024484,0.00667549817003898,0.00494615932505948,0.000731649393775236,-0.0106073005763221,0.0209214068111252,0.013777356550581
"1803",0.0140557154983383,0.0202833334839578,0.0255732478603772,0.0170190045174796,-0.0150420685404985,-0.00768412309214161,0.0122806799248603,0.0160818578278172,-0.0123570503223529,-0.00377495795619198
"1804",0.000906057002560745,0.00124229505203122,-0.0111780009982948,0.000760852455685468,0.00214210568880047,0.00107829537526416,-0.00129979668126345,-0.00311750086318274,0.00163200195387003,-0.00833649397690217
"1805",0.00229026261434839,0.00868675015879905,0.0191303369968148,0.0141878573764207,-0.00984972647891424,-0.00430803686667924,-0.00477210544743012,0.00793842742354545,0.00993094118962645,0.00917079873772564
"1806",0.000425118485881226,-0.00676659006653391,-0.00682606536155794,-0.0127402874701181,-0.00628777676870906,-0.00432711047709944,-0.0113340788181938,-0.00119354764487245,-0.00829685808245906,-0.00454367128187516
"1807",-0.00053094345692839,-0.00639953168050045,-0.00429549111239536,-0.00683215006325766,0.00141687555639836,0.00108599260823383,-0.00367412410706247,-0.00931915098388647,0.000309931065455959,-0.00836828159099012
"1808",-0.00494286090015428,-0.00498640287619689,-0.0103537912131164,-0.0112097397347292,0.00264022254694218,0.000987509757696348,0.00545804991517596,-0.00651217015991012,0.00565318649217117,0.000383577422433889
"1809",0.000267206451574964,-0.00292364823562663,-0.0095902246874221,0.0020609064135837,0.00696017904490231,0.00394212574718433,0.00220070931627281,-0.00534090572942103,0.0146310949127437,-0.00268401243046767
"1810",-0.0112132929063483,-0.0215704426655455,-0.0167252778768339,-0.0179993773157696,0.0134506177942306,0.00589043636339071,-0.00322077423173772,-0.0126921934530783,0.0034153917507358,-0.00461366569400934
"1811",-0.00280803334075752,0.000856165778564622,-0.0116383322058891,0.00549857413868993,0.000184325415711006,0.0000975194938450663,0.000293690768563337,0.000741278331982009,0.00673170677617474,0.00540753876743816
"1812",0.00904351995052721,0.0130452816106914,0.0108697050244639,0.0122396914034009,-0.00746411145822201,-0.00400120131594184,0.00161511622361554,0.00914059055659777,-0.0109692481907178,-0.0111410364454776
"1813",0.00713792085091214,0.00865523060200002,-0.00089610802049056,0.0138923880792252,0.00362052897857756,0.00244911767457157,0.00439732292982153,0.00538542700150724,-0.00774843518496227,0.00505051615747321
"1814",-0.00532869707489236,-0.0146503801211147,-0.00538137120078896,-0.0213141909676499,-0.0077702189682799,-0.00928558487564135,-0.0176590769628013,-0.011200226609252,-0.019369155541615,-0.000386463282109228
"1815",0.00583946808480129,0.00127432590810672,-0.0144270835348299,0.00440747593938617,-0.00177111120231654,0.000198183185299294,0.00133714237516447,-0.0123125040597395,-0.00179557348100801,-0.00464046671164819
"1816",-0.0038785086937525,-0.00318196523071534,-0.00457482376311025,0.00619514032981439,0.0108336884158178,0.00187359108158103,0.00816027122455698,0.00170640105365072,0.0047708430723381,0.000777070152832904
"1817",-0.00413541803792317,0.000212965877965265,0.00367657740440541,0.00974866689127452,0.00711429204953262,0.000394187090041909,-0.00588635115522118,0.00325668833618198,-0.0178251808373535,-0.000388273345873769
"1818",0.00474573307582493,0.0129786659641644,0.00457881107816926,0.0114330887844514,-0.0037617418846001,-0.000590969669736152,0.00732241006587686,0.0099875607420099,0.0018228245363765,0.00660197167429399
"1819",-0.00719199570626683,-0.00189041290164804,0.00729265029123094,0.00226073550359507,0.00782831848852905,0.00423459531647796,-0.0111494811449834,-0.00494455323488718,-0.00791076630295806,-0.000771634106060737
"1820",-0.00210844912493469,0.00273564383262914,0.0144796049567577,0.0130322759317878,0.00502541518488808,0.00098039565005581,0.0048107242064932,0.00993793443923807,-0.0065386171265891,0.00888022757835838
"1821",0.00492970734044684,0.00629599427149552,0.0107045680267512,0.00791706389937574,-0.00563726701589229,-0.00352647759073943,0.00658291314980408,0.00984000633684512,-0.000240773745590395,0.000382775466384988
"1822",0.00819444866590624,0.00688202865498511,0,0.0066272722609666,-0.00246824062817985,0.0000986629555923546,0.00579665081519742,0.00292342431103254,-0.00762682253736069,-0.000765021771425012
"1823",0.00663089712076403,0.00683536546619412,0.00264781679101378,0.0117042812608164,-0.00854645785044184,-0.00206860206648352,0.00635440415298305,0.00218604992530369,-0.00177980744454487,-0.0122512563764504
"1824",0.00334661103921841,0.000411239730689683,0.00880292659285509,0.00192842317635944,-0.00574672404647758,-0.00434228016879812,0.000146778059942676,0.00799799845295013,0.00753708572442724,-0.00232554975998711
"1825",-0.00132332984693917,-0.00267327633073688,-0.00523560879658203,-0.00384898037654124,0.0043815457910501,0.000693689355305782,-0.00352360545174835,-0.00384710978440939,-0.00321751930501923,0.00815851687320612
"1826",-0.0118225318070967,-0.003711246931284,-0.0043859462756668,-0.00265649911188492,0.00668297877607826,0.00614163714350346,0.00397818980935849,-0.000724076720451383,0.0133150583168988,0.00462429368806183
"1827",-0.0110512645514143,-0.00393217560970338,-0.00969161785873429,0.00435834926303369,0.00599281709798705,0.00236232933433822,0.00102723318258224,0.00458936697043333,-0.00525600063709475,-0.00230146453460378
"1828",0.00412278076571293,0.00332443595240139,-0.0213522907317479,0.0115718860744736,0.00238290260308927,0.001375305777779,0.00557113150055866,0.00264467814297542,0.00944673734859536,0.0115339861699637
"1829",0.0107508467289514,0.0132532574150801,0.0145454976441539,0.00762641267437636,-0.0049372719431231,-0.000294463510875809,-0.000729090129865773,0.0115111211565668,0.00182412568242118,0.00266054900521828
"1830",-0.0210058302411522,-0.0183937266986323,-0.0286738444599149,-0.0106433999144944,0.00928083046173334,0.00421853191803789,-0.00889991637331677,-0.0113801231798667,0.0054623337555415,0.000379147925316126
"1831",-0.00900860444802953,-0.00666248867503216,-0.00369004132898365,0,0.00810248948804815,0.00205151249085422,-0.00603547552435713,-0.00167836125132892,-0.000629887400521389,-0.00454719271475734
"1832",0.00787820466911504,0.00482092697607417,0.0138888799896597,-0.00215153611964058,-0.00261898787488479,-0.00155971544297395,0.00370243353986766,0.00384354705405276,0.00724807374143221,0.00913592825592224
"1833",0.00688768675426354,-0.00438060835310661,-0.000913293674612681,-0.0150933642271043,0.00624752171756304,0.00117159741770645,0.0106242232940819,0,-0.0184591320838347,0.000754344303005805
"1834",0.0104779025063215,0.0111041712519608,0.0191956367156165,0.0126490879079495,0.00125998179627618,-0.00156048917962104,0.00598614549709087,0.00885363653552962,0.000398462035197555,0.0018846720080643
"1835",0.00139653289671138,0.00580189074532478,0.00269046217307145,0.0091277174310922,-0.0109643143888561,-0.00566573995114072,-0.00275761491193049,0.00450656969896723,-0.00629282295449407,0.00225738301863121
"1836",0.00348735023188507,0.00185409417460147,0,-0.00618880522246545,-0.000818047182561843,-0.000196644323885775,0.00422072697246301,-0.0028336848087227,-0.00408819238476954,-0.00337844807662935
"1837",0.00454452942432582,0.00658031134429859,-0.00715557053068494,-0.00263464492235699,0.00336508950720571,-0.000392755391060873,0.00333309073269406,0.00497291645215991,-0.00370250327917743,-0.000376565178978328
"1838",-0.00234189295688825,-0.00326864695749451,0.00270275608154424,-0.0072048783926123,0.00571003842985696,0.00255559571862252,-0.00303303416583101,-0.00282734659238848,-0.000161552756192895,-0.000753569186683123
"1839",0.00202719022640729,0.00143467311444878,-0.00359409381426457,0.000967640598329211,0.00189267315676211,-0.000293778789080656,0.00333225291545558,0.00307173414320649,0.00646409168610051,0.00603313866066468
"1840",-0.00819869412694174,-0.00450256953711037,-0.00631167744941097,-0.0135331776206667,0.00143929100457574,0.00137289608824509,-0.00346574573708769,-0.00494701129744535,0.00698460191047867,-0.00412292080413723
"1841",0.00316711924311419,0.00328928034149212,0.00544437595293412,0.0048998925788879,-0.00485049569799589,-0.00146903744987026,0.00521673502472941,0.00378784297637869,-0.00438493980706378,-0.00338731004097692
"1842",0.00465529200222203,0.00840170425955433,0.00270773490793852,0.00950740510783987,-0.0013538796378173,0.000882723650467376,0.000576655449463281,0.00589618323064234,-0.000160121720694795,0.00264346846756669
"1843",0.00298282840740227,0.00792525701684754,-0.0027004228786438,-0.0019318150415617,0.00415810200349243,0.00264565824801455,0.00446619420907557,0.00140699096014196,-0.00512574078867745,-0.00527299793137248
"1844",0.000106066884610456,0.00201622996422635,0.0126356215771399,0.00120957874614191,0.0107276492449297,0.00287947857829152,0.00774525973781914,0,-0.00338108192415798,-0.00757290238187724
"1845",-0.00143361832127853,-0.00321932113936674,-0.00178273062415291,0.00555826292791006,0.00615942176887452,0.00146476445827926,-0.000426941076854925,-0.000234016452356878,0.010177665343029,0.00267073913185523
"1846",0.00191423135011459,-0.000202003759240732,-0.00267852564066917,-0.00552753941052186,-0.00603312162284841,-0.000585042227234545,0.00355963819034799,-0.00117127176248477,0.0092755718739097,-0.00228319130765142
"1847",-0.00870384758998577,-0.00222073381798493,-0.00268574418977974,0.00459175230557607,0.00401697441663118,0.00117069238983936,-0.00368897732891948,0.00422054727351795,-0.00190142606638066,0.000762844652970829
"1848",0.00588934291238363,0.00364215826801639,-0.00448848522562539,0.00529241026674754,-0.00355630166240106,0.000779801731829899,0.0116776560433074,0.00817183361863894,-0.0143673992451008,0.00266768573702603
"1849",-0.00106461430707472,0.000806647897340085,-0.00360658368689615,-0.0023930789940636,-0.00428269714541885,0.00107089366343049,0.000563241961169858,0.00115779908357183,0,-0.00304070567216974
"1850",0.00149197341670182,-0.00423051447761758,0.00814468071973828,-0.00167911300063317,-0.00322603674812838,-0.000778360573503667,-0.000140766825680871,0.00277577564208276,-0.000563743264294869,-0.00495612882897922
"1851",0.0097359921931004,0.00809226452699474,0.000897716923160319,0.0168189295040717,-0.00404516723273274,-0.00262843831480397,0.00211048222968291,0.00553631292060053,0.00676876723237352,0.00229889807629657
"1852",0.000895953975583286,-0.00220755749566026,0.0134529314968104,0.00378065956663143,0.00866511736298126,0.0039046034797352,-0.00589717496673881,0.00206500692409173,-0.00272133819879405,0.00458713250180853
"1853",-0.00473798074657072,-0.00140803225802921,-0.00530976551228146,0.00706222027424941,0.010827872275315,0.00456877110291765,0.00254248360558362,0.00251826289632739,0.00971107559728845,0.00456614763446561
"1854",-0.00878020309320837,-0.00382664829118773,-0.00978646453317766,-0.00935047517217258,0.00796739103349253,0.0035811190384738,-0.00169072616874344,-0.00159867070798481,-0.00826644159075485,-0.0060605625859117
"1855",0.00346836615872781,0.00141514081452421,0.0017969474276609,0.0132140399846488,-0.002810878863446,-0.00212164507308099,0.00733845957486978,0.0036596817870469,-0.00216395773416589,0.00114331630053921
"1856",0.003669258422623,-0.00141314102098866,0.00179364972380047,0,-0.00739791733506112,-0.0012561276462999,-0.00364241082371053,-0.000227967682430719,0.000642586345381391,-0.000761353473580639
"1857",-0.00630483450229335,-0.00545891680774468,-0.0116383322058891,-0.00815108655977592,0.00221832535455113,0.00290262180355905,-0.00309343839909548,-0.0093459098081653,0.000882966754166548,0.00190477512353748
"1858",0.00842437349455061,0.00833489336748006,0.0117753779665133,0.00774845242120059,-0.00610870683646825,-0.00154344162970887,-0.00394922954528654,0.0043720889287,-0.0024059908187346,0.00190111471928089
"1859",0.00243223553199323,-0.00100811498211328,0.00984779477801911,0.00698992826197475,-0.00142534567578545,-0.00106298048788434,-0.000849547147671936,0.000916291622828469,0.0022509767847172,0.000759081054928057
"1860",0.00400861545121312,-0.000403633412779714,0.00975185958931957,-0.00185112559559208,0.00535220742408127,0.00203142234885734,0.00751112328477266,0.00595095456184991,-0.0012833560805865,0.00227528168495428
"1861",0.00614667227702848,0.00868167135896214,0.00790162931902283,-0.00857674376296846,0.00585628702203134,0.000289694176745403,0.00604868858730345,0.00227531542174408,-0.0213637776666328,-0.00832387743504726
"1862",-0.000731168860092168,-0.00460373922302382,-0.00435535803942266,0.00584523889969679,0.0123499534708813,0.00550050573239735,-0.00405503693546805,-0.00567520094380325,-0.0053344358692563,0.000381450015833007
"1863",0.00517290156373962,0.00361964915605628,0.0113734712643345,0.00278939707238424,-0.00531509088038173,-0.0012475786594206,0.00126361240527495,0.00525082459263859,-0.00214517332042496,0.000381422326485303
"1864",0.00161142125669156,0.00140255109695331,0.00173020190525741,-0.0136764667108661,-0.00043848502137489,-0.000768837274531475,0.004907334118748,0.00272584925121921,-0.00421698355850864,-0.00762479245482162
"1865",0.00114183694175263,-0.000800224739854416,0.0120897772377941,0.00305527989704091,-0.0074335919765921,-0.00457607621506906,0.00181441069246757,0.00385042113605616,-0.00606163746574784,-0.00115257963929916
"1866",-0.000518316134909713,-0.00300382673429755,-0.00170641596436916,0.00562320942578176,-0.0123047813327823,-0.00503235779784583,-0.0012537036498258,-0.000676861277936425,0.00258984968896869,-0.000769141123897699
"1867",0.00202282124909114,-0.000803278521829598,0.00683754411289228,-0.00559176575587639,-0.000269474049539586,-0.000778134801900587,0.000976146500597519,-0.00293529386561886,-0.00208315970197215,-0.00269442259198116
"1868",0.0065218897176591,0.00824114697798173,0.00254676302809909,0.0105436220917847,0.00044853861936911,0.00146016633578405,0.015603271728067,0.0040759455279189,0.00751504663468516,0.00115791773421514
"1869",0.00478273409338992,0.00737645650652752,0,0.00996979353856009,0,-0.000777616277002013,-0.00205769409270651,0.00902117849876727,-0.00041441238473694,0.00424041755856797
"1870",0.00102401499422156,-0.00178117093372754,-0.000846787938743487,0.00367303770446425,-0.00143379588869919,-0.00145890919969083,-0.0107217520145395,-0.00447005935350731,0.000331655747187964,0.00422274939862954
"1871",0.000102205537759081,-0.000792926957389417,-0.00847453989177105,0.00526084991600584,-0.00367982121191801,-0.00175382795225487,-0.00514080164797626,-0.00202102427028594,0.00613341887884933,-0.00267588302880972
"1872",-0.00347674757834726,-0.00674611466738284,0.00256398736658481,-0.00341304385769714,0.00180184551664797,0.00136637511961935,-0.0040504172322583,-0.00517372854534892,0.000164799408228111,-0.00268298369309872
"1873",-0.00707968880237941,0.000199712355313242,0.00341015857336502,-0.0047945153863389,0.00890118306005361,0.00389826810628269,-0.00294483072466423,-0.0027140407520081,0.0101309196892869,0.0142198340612605
"1874",0.00304839098259535,-0.00139799693801768,0.00509764171367055,0.000458952254876133,-0.00053470266655764,-0.00194164727948398,0.00253141778650834,-0.00385513565577,0.00260926290451113,0
"1875",0.000824126259973079,0.000199855345329514,0,-0.00458630951745187,0.00249669705386446,0,-0.00505053104888986,-0.00455267149096272,-0.00439168025692638,0.00303140980953276
"1876",0.00277972057038323,0.000200008702963883,-0.0016905256577805,0.000230440916557217,-0.00791626988090322,-0.00418267714245324,0.00112839027103062,0.00114352494525938,-0.00114359583636003,0.00113334305133139
"1877",0.0073394977473189,0.00799679161103506,0.0135476929417415,0.0110547484697605,0.00771035998617009,0.00527477922226782,0.00619701295435959,0.00776599061653838,0.00318939322202638,0.00415104216286699
"1878",0.00112100840342944,0.00238020398817884,0.0175438831794341,-0.00569449302324077,-0.0128115138651992,-0.00252593959077607,0.00769869981540494,0.0031732692284443,0.0348088698917237,0.00977074474588324
"1879",0.00203020821444189,-0.00257227202172317,0.000820996418668285,-0.00206203744328226,0.00757057809758854,0.00116840272064223,0.00347282412393901,0.00247021474684139,-0.00346622020692899,0.00186078579704874
"1880",-0.000306100033490964,-0.00178541098273921,-0.00820341102293665,-0.00206600780209631,-0.00313089621401985,-0.000681335121090476,-0.00235317389570466,-0.00547574519332217,0.00276678260869567,-0.0037147358734172
"1881",-0.00602428716892045,-0.00765390411662836,0,-0.000460219141565799,0.0101393608547271,0.00408948260403008,0.000461829224696064,-0.00183517144763723,0.00102487191209888,0.00149140393515124
"1882",0.00451985452743853,-0.00123377489941867,0.00349779746938728,0.0021111008057848,0.00257594881410039,0.000969694167155755,0,0.00666501669400565,0.0000787131813189124,0.00148918296182177
"1883",-0.000715657935823621,-0.00144150114204644,-0.00331962431161426,0.00115722382817163,0.00478426639796803,0.00261522018888916,-0.00111910214926259,0.00616444477671907,-0.00204736596657007,-0.00408908711055656
"1884",0.00194413675936977,0.00123727633734183,-0.00249796490817478,0.0023119570982908,-0.00149907853422093,0,0.0060207669025627,0.00476504732637251,-0.000552347497379868,-0.00186641921430597
"1885",-0.000510710356701805,0.000411931947262412,0.00500853251993716,-0.002767917551876,0.00247290131615707,0.000773523992263936,-0.00083500243889445,-0.000902991409806653,0.0108952230887345,-0.00598361722093199
"1886",0.00669322735312194,0.00885316863938268,0.0174417946175502,0.00948403969185341,-0.00837294078905415,-0.00326959713553565,0.00250711822897887,0.00565069902597792,-0.00265538908612728,-0.00300977948909364
"1887",0.00101497009873142,0.00102031226957733,-0.00244886790916554,0.00595774561970175,-0.0106872779388185,-0.00407576132860543,-0.00111134092134824,0,0,-0.00188676673158761
"1888",0.00491828082568579,0.00550445415636047,-0.00327353274621645,0.00592269503313836,-0.00360125467622652,-0.00204571690477851,-0.00472962317366654,-0.00134858969476326,-0.0042286062074065,-0.00189041117318534
"1889",-0.00348155191122101,-0.0115570244773275,-0.00738914232481003,-0.000679235025344505,0.00731846383979406,0.00244090927653051,0.000978525948034825,-0.00472615854899971,-0.00110103016354102,-0.00795447621105305
"1890",-0.00642997539736823,-0.0133333362293296,-0.00330839155671014,-0.00453232836029371,0.0112120165712069,0.00457800660064156,0.00307154251449226,-0.00904615482896631,0.000393662424665209,-0.00267273931650935
"1891",0.00448420653444015,0.00395017330606029,0.00663883794805598,0.00569103602539234,0.0007985512351949,0.000193344737687617,0.00222714052994588,0.00890023940548268,0.00605962068151422,-0.00689125536772417
"1892",-0.00395667374330066,-0.0124248858487093,-0.0173124768946333,-0.00543242753358364,0.000265398789426552,0.0021327751870992,0.00319467132719087,0.000678752549222006,0.00547557119760866,0.00154199887714679
"1893",0.0013752485508991,-0.000629126903002875,0.0016779144595751,-0.00113770919211942,0.00637955195279227,0.00164409402052956,0.000692183216005615,-0.000451966127483439,0.00186716985428803,-0.00885304054897218
"1894",0.00503515236972629,0.00692398723871923,0.011725404094322,0.00774674742316717,-0.00431408233515507,-0.00222095656717314,0.00456551308705366,0.00407047022237705,-0.02376143829602,0.00388352215418641
"1895",-0.00187258925057376,-0.00416748681207413,0.00331110718196048,-0.000678546869511854,-0.00203380292125521,-0.000871026649221562,-0.000275334464242549,-0.00045046167350915,-0.00946549467494828,-0.00928428552675742
"1896",0.00370145877032368,0.00795129813276474,0.00165015801680157,0.00248877379853663,0.00531621274500416,0.00145314357631565,0.00371933530467006,0.00743562534759445,0.00353330124093221,0.00156178810632168
"1897",-0.0113663163721089,-0.0153621856135829,-0.00658978057148729,-0.0187317542580737,0.0126037699041992,0.00580378135211523,-0.00590151488316404,-0.00849912184379198,0.0169640312317834,0.00233922971859379
"1898",0.0102195009052439,0.0078011306143857,0.00497512607933115,0.0156394379207951,-0.00322081556606579,-0.00201931845746084,0.0088359581899784,0.00924851782663927,-0.00755369447017684,-0.00661216291621969
"1899",-0.00187127861403558,-0.00460264382323583,-0.00165004459920248,0.00339676942829992,0.00497760065517849,0.00028866792201887,-0.00287401400390042,-0.00223513118886354,0.00166494097355763,0.00469848805988504
"1900",0.00435787180444458,0.00483397980996947,0.00330565709764485,0.00925295580890451,0.00208555214707218,0.00125271294385199,0.00425464257067554,0.00403239088171237,-0.00474907407785574,-0.00428688944394529
"1901",0.00221984521217489,0.00104590497430523,0.000823866940642848,0.00089450148860748,-0.00130112709607666,-0.0000965106147188255,0.00218705271446229,0.00401570360614412,-0.000954310497126021,0.00273980957205633
"1902",0.0000505509461088405,0.00522347103018928,-0.00493836312063745,0.00446812796145402,-0.00746601584430862,-0.00404163960176174,-0.00259119223912907,-0.00177754724656864,-0.010109894679751,-0.00117094414663099
"1903",-0.00468152100199115,-0.00706706107611987,0.00330848251593219,-0.00400347809852941,0.0118085654748776,0.00386519466693858,-0.00560544512977301,-0.00823682804401638,0.011580241440776,0.00390772288067054
"1904",0.000404224561015631,-0.00167465698002334,0.00577089362600236,0.00692267125849066,-0.00138318588233188,-0.00115504398697708,0.00604932892009358,0.00157133884875305,-0.00166944111877387,-0.0019462560111887
"1905",-0.00429723596770482,-0.00293559661790144,-0.00245915223010207,-0.00598801713304442,0.00363590838196504,0.00134870535633458,-0.00464630384507447,-0.0011203855389984,-0.00302599931476344,-0.00312016237850077
"1906",0.000152443164238125,-0.00210297535073878,0.000821768309770432,-0.00490851452865859,-0.0138872297799564,-0.00702465259151031,-0.00096131067779448,-0.000224433664764989,-0.00295523170020529,-0.00430358089483418
"1907",-0.0197481944243147,-0.0195996925583148,-0.0147783749367313,-0.0174888543341852,-0.00297446710421001,-0.000290704379270146,-0.0144312073306559,-0.0130166387191458,-0.0115357123842711,-0.0051080660694437
"1908",-0.00305548871729289,-0.00795362997936455,-0.000833066351322298,0.00547716220299543,0.00774099427755925,0.00588588567260517,-0.00195226555010664,-0.00250079301392514,0.0080233244835346,-0.00789890821798944
"1909",0.00722064254245214,0.00476689651937434,0.00166786580085643,0.00930553510705057,-0.00261862978002769,0.000578846170027569,0.00600807853368357,0.00364713680251461,-0.0031355443753549,0.00756371398691158
"1910",-0.00969614130042251,-0.0116450534193068,-0.0158201849839582,-0.0152913438712744,0.00323807354033656,0.00048239218730517,-0.00888846934628462,-0.00885766355420681,-0.000967779675260627,-0.00474118489242559
"1911",0.0003125418890495,-0.00218228477643168,-0.00507616704416425,-0.00685096650880934,0.000610985194516633,0.000868906310670825,0.00182139206981669,-0.00779108774231496,0.0145313228094457,0.00635168079479187
"1912",-0.00541468747784324,-0.0113711042281501,-0.00340129939586553,-0.00390880321496889,0.00932813977833669,0.00452895562751454,0.00153869587675026,-0.00461889534193827,0.00405826377111906,0.00197235968110299
"1913",0.0115687431019533,0.00906897976885679,0.00170664152001221,0.00900261829840865,-0.00215906775463559,-0.000863506215697529,0.00754198036239995,0.00556839424054556,0.0000792677127912089,-0.00472426408615978
"1914",0.00289792853911774,0.00197265917897571,0.0093694355803764,0.0128119981679358,-0.0000864593999022611,-0.000480231217428462,0.00554480926411993,0.0108447601937882,-0.00182267213213938,0.00158217528215698
"1915",-0.00139291731385294,-0.000437396983988925,-0.00168764060433313,0.00112915079807885,-0.00649316234796737,-0.00144121346454473,-0.00289501214091747,-0.000685075689544901,0.00023816291075085,-0.00631915096339819
"1916",0.00676869831348492,0.00415832562626894,0.00845314169727529,0.00541526804102843,0.00653559905366397,0.00327093742416196,0.0124430273449663,0.00799487833767776,0.00166679104161904,-0.000794901731337117
"1917",0.00472188399874462,0.00566701491501664,0.00167641553019027,0.00157085112429023,0.00805112930960439,0.00201400818181763,-0.000273260328101821,0.00702440655821746,0.000871640274286101,-0.011933134359741
"1918",-0.000204312108424531,-0.00130039542230431,0.00167354084598714,-0.00268871163227069,0.0109068978254405,0.00401861079816679,0.000955995615397054,0.0036001407279771,-0.00657109502923114,0.00402575128422056
"1919",0.0083795366896442,0.00781240425631013,0.00334171925042837,0.00966062478763763,-0.00993989653234484,-0.00314502221855306,0.00927977200472929,0.00470870217038155,-0.00414411848555662,-0.00842021728674447
"1920",0.00521875955105222,0.00193820793376021,0.000832716012798995,0.00467293445181172,-0.00308918046411555,-0.00105132648656758,0.000811180664066713,0.00490986589568609,-0.00224070904481988,0.00202189146360765
"1921",0.00267154096279776,-0.004298352892249,-0.00582363615512493,-0.0019931510673098,-0.00163504094103029,-0.00296736535762587,0.00486347811046683,-0.00621832472781969,-0.00368943695861412,0.00282482003879458
"1922",0.00291579851013934,0.00561176772625993,0.00502085260007701,-0.00421695465151795,0.00560414406811116,0.00211211015725721,-0.000941092723526382,0.00335216352851986,-0.0107873449461653,0.00241449533829319
"1923",-0.00155411699100905,-0.0051513919285836,-0.00749382605069093,-0.00267405102684037,0.0055725355727525,0.0000954192885884719,-0.00672864244907168,-0.00178175124713997,0.00252282721002994,-0.00160580016755862
"1924",0.00507050333028092,0.0101404282470239,0.0033559211756149,0.00737414751104959,0.00375125544891342,0.000766773010544064,-0.00040645716645038,0.00401570360614412,-0.00365292631458847,0.00160838290910359
"1925",0.00064949981623208,0.00170863652604392,-0.00501681508627738,0.00598934532265494,-0.00322748028819253,-0.000191490021558827,0,-0.00133275429430091,0.00496985505898406,0.000401439712543361
"1926",-0.000399212187565778,0.00405131881211473,-0.0042018125916361,0.00507181275016189,0.00852081613077682,0.00277599898410741,0.00162638773023627,0.00311515828026709,-0.000243194166894112,0.00160511449347278
"1927",-0.000549647024469135,-0.00594615070700566,-0.00253160010866116,-0.00987276341619825,0.00523945425465655,0.00133645077981459,-0.00094681499733773,-0.00510232150350287,0.00551410963347387,0.000801271114856617
"1928",0.00284836742417083,-0.000213710013883706,-0.00169201691598242,-0.00155103615637342,0.000672346906914756,0.0000955311819754723,0.00501136848606687,-0.00267549923302568,-0.00112902419354843,0.00200165638693472
"1929",-0.000498526733105797,-0.00085484681047121,0.0101694246306123,-0.00155359754527995,-0.0172506921569212,-0.00638865499908337,0.000538733565223382,-0.00268276924397703,-0.0178427174403138,-0.0143828316073027
"1930",-0.000548401524546049,0.00940980024381388,0.000839095614485252,0.0131141137159305,0.00556862425101579,0.00144155933623513,0.000269813254244466,0.0100872768968747,0.00411015200805331,0.00405353459188329
"1931",-0.00144619665827983,-0.00508471724588666,-0.00335301541861688,-0.00263289712988135,-0.0121827188329975,-0.00355078150406574,-0.00188542931735136,-0.00754550270816667,-0.00548505107678998,-0.00403716978450852
"1932",0.00449517896625129,0.00212957262662661,-0.00420534682122364,0.00857892731857457,-0.00189747161513876,0.00028868551105532,0.00944426034679213,0.00178913924068813,0.00477440719193911,-0.0016213804612808
"1933",-0.00258547886093663,-0.0131747825434131,-0.000844393734122373,-0.0117774230304565,0.000432276557848832,-0.00105893752520869,-0.00173768326036816,-0.0111606255613018,-0.0108962397328566,-0.00487208260272087
"1934",-0.00633133349893944,-0.000645756861875957,-0.0084531416972754,-0.0123591981359261,-0.000777572082963029,-0.00231295936916309,-0.0053553192630228,-0.00835226040537485,0.00115961232933959,-0.00815990734283745
"1935",0.00376263120480225,0.00409381353290428,0.0110827051364992,-0.00424591214682601,-0.00631004590124318,-0.0025125056587002,-0.0138645008228787,0.000455249813114733,-0.0050467525842619,-0.00699312305008326
"1936",0.00114978909332941,-0.00450636775998392,-0.00252946534234466,-0.00673247883477579,-0.00330560930244184,-0.00125863092498679,0.00122837147629085,-0.00750859611322197,-0.00656910848878922,-0.0049708498179174
"1937",-0.00584155690409227,-0.000646833171491834,-0.00338119625600142,-0.0106190933566749,-0.0104728497830162,-0.00378213873297673,-0.0287662282558661,-0.00320955475768003,-0.00912366276786081,-0.00791018072039307
"1938",-0.000753246755016757,0.000431365877238354,0.000848091097809256,-0.00502396914538783,0.00149963287351063,0.00184948130263485,-0.00407097503011566,-0.00850924029643496,0.00219633389583551,0.00125898658360835
"1939",0.00753846956190918,0.00366538411917672,0.0016948846895477,0.0130823715779553,-0.0040513627290657,-0.00029132509391383,0.0074704186875767,-0.00139220700037079,0.00160150877951359,0.00922045596687138
"1940",0.001346934027882,-0.00386690184506566,-0.00846020087612909,-0.00928859309820562,-0.0025642828648037,-0.00252706946769499,-0.000699656543412308,-0.00627161514852337,-0.0108558527163871,-0.00415285260395082
"1941",0.00532995673854808,0.00927340766156148,0.0059727761660382,0.00137203672670583,0.00319160829538645,-0.000681926576165837,-0.00727983636317331,0.00467478008265809,0.0020418410580072,-0.00959132395730922
"1942",-0.000901115515094308,-0.00491444530723795,0.0016963454245893,-0.00753594068931895,0.0127248682634813,0.0038023750561873,0.000563870708063297,-0.00503663256407916,-0.00585840555152328,-0.00294732818754173
"1943",-0.00772302006886816,-0.00365053021373896,-0.000846817831226754,-0.0151862983648804,0.00122196692274956,0.00213718272594732,-0.00887921261037228,-0.00329635082906143,-0.00204968834399821,-0.00844604763001489
"1944",-0.00572420605636192,-0.0129310117501775,-0.00169490798821303,-0.0056075848213355,0.00618774718726089,0.00213188694676525,-0.00568833623435927,-0.00685113531231718,0.00641848534734257,0
"1945",0.00782793806337589,0.0045849019230535,0.00594219117938,0.0143326240232131,-0.00554313941744766,-0.00280476398467966,-0.0010102919647057,0.00404410485261297,-0.00467682831083038,0.00425901741067269
"1946",-0.0161354098987053,-0.0163006321820667,-0.00253160010866116,-0.0217744587825885,0.0118454901552443,0.00484995413006817,-0.00491186153604795,-0.0156363340030403,0.00290470731555637,-0.00212041208275215
"1947",0.00794542957868405,0.00419804115327538,0.00761419241813788,0.00449925359648451,-0.0014633881816859,-0.00212369779055144,0.0110336700771267,0.00890469953768691,-0.00281115088858641,-0.0016999779678657
"1948",-0.00181913508414688,-0.0074807701387547,-0.00587751600135389,-0.0202732209907432,0.0080173383437423,0.00319223416307901,-0.000287204124269635,-0.0102574517752779,-0.000256270293119143,0.00595994531177846
"1949",-0.00263229852684543,-0.000664874229936108,-0.00591198679657512,0,-0.00564424192856716,-0.000867814435637659,-0.006032554972769,-0.00192816320094313,-0.00700675046575028,-0.017350806458111
"1950",-0.0135520664973633,-0.0126443295012667,-0.0161426778798385,-0.0204524918930185,0.0193908295856313,0.00840187882938337,0.000577934675108471,-0.0074863603545936,0.00481884523551201,-0.0034453030602557
"1951",0.000154377630292801,-0.011233353412135,-0.0189984510465246,0.00540418000950349,-0.00871183977908974,-0.00297240391008435,-0.00158862234230872,-0.0065687487146977,-0.000256906746345154,-0.00388940490539325
"1952",0.0110095250487725,-0.00431719572827094,0.0123241340750511,0.00855094439142912,0.0042662323859568,-0.000288543186848123,0.00679853071590886,-0.000734895702450444,-0.0182456487621321,-0.00954442786635024
"1953",-0.00117088012570765,0.00821543290952187,-0.00260893525720995,0.0130816022615972,0.000594528156440344,0.0016352955597172,0.00129325080004628,0.00171557006073741,0.0123898262595776,0.0127025911314935
"1954",-0.0154360882313302,-0.0212765923451498,-0.0061027919148865,-0.00884757247757073,0.0135010779708988,0.00585846625139963,-0.00588308549137939,-0.00831928317760122,0.00284410930659407,-0.00389276939652727
"1955",0.0174891914958408,0.01919507159281,0.00614026467248507,0.0149576468867214,0.000251306576564359,0.00353188883713296,0.0190531422995122,0.0148039425174482,0.00953936052303739,-0.00390789288984161
"1956",-0.0198329243540586,-0.0297253947830579,-0.0252832553106828,-0.0156878424245721,-0.00435544909183105,-0.00171239746139151,-0.00127505571929554,-0.0133724119867671,0.00144716096495134,-0.011769807888793
"1957",-0.0114143630265635,-0.0137981588129297,-0.0143110620498899,-0.0217341273773347,0.00992710306843692,0.0039074301820321,-0.00141789658928393,-0.0056674062365234,-0.000425051006673338,-0.00352893522585584
"1958",-0.0164269413749547,-0.000236889983532107,-0.00907456944861107,0.0101209218541483,0.00608053740760583,0.00522123820007869,-0.00170436157986331,-0.00322160553782214,0.0079088445585116,0
"1959",0.00154734296838122,0.00071161969677136,0.00641006532925248,0.00586521736899637,0.00654072079777834,0.00198323362545927,0.0150803105661357,0.00273464545452806,0.00059060919483489,-0.0150509295657192
"1960",-0.00676630924535204,-0.0106659518999835,-0.00545913609228244,-0.0126337920219065,0.00789681431775935,0.00565494055202276,-0.00700793421636658,-0.00223161318867771,0.00337298265867214,-0.0125843292251807
"1961",-0.000857928905226957,-0.0103019420536546,-0.00365981206604338,-0.00910413143206201,-0.00636582203519143,-0.00271783626397126,0.00268203532976274,0.00447283437968071,0.00193296078549388,0.0100137531760711
"1962",0.0118106472997039,0.0220284865255622,0.00459141157870846,0.0111744733723367,-0.00558525369115048,-0.00291322341847466,0.00506744333579778,0.00890698673417778,-0.00192923165635606,0.00360527101475738
"1963",0.00970968798236838,0.00450012052003368,0.0201097776978749,0.00294699830539269,0.00363427209989831,0.00141368773699524,0.0142856734867693,0.00882774805958952,0.00680733686540624,-0.00718459324177123
"1964",0.019811125614875,0.015090779030706,-0.00179218065299225,0.00416254683504325,-0.00798287969936684,-0.00272926287255704,0.00952782034571631,0.0109380428085741,0.00183634386052556,0.00814114085177753
"1965",-0.00711075743253153,-0.0111500092001915,0.000897649807543033,-0.00658353026180203,0.00107814674548545,-0.000283168050011939,-0.000410137819130574,-0.00769407593866367,-0.00566573085316779,-0.011215776547182
"1966",0.0116246307706724,0.0136249451133041,0.00627803656955805,-0.000245632956918262,-0.00886678301234689,-0.00415355868459288,0.00752604425463343,0.00993458443744522,-0.00687111636906701,0.0117966179513764
"1967",0.0076952393446279,0.00463504936876435,0.00356502233636835,0.00712028729700065,0.00100306461518573,0.000852992311288325,0.000407443827152409,0.00239912656490371,-0.00143434866944858,-0.00627794142929505
"1968",-0.00137442829706447,-0.00553632720278618,0.00177606917816542,-0.00780128752162867,0.00183806966592415,0.0010420516457994,0.00597298134585267,0.00191468139568474,-0.00245035914576019,-0.00270768346460881
"1969",0.0114700444078752,0.0153097614295479,0.00531934599219874,0.0201474590394126,-0.00625327098855122,-0.00246006443966029,0.00323892765950795,0.0102728089519206,0.000338810779922261,0.0081448253341041
"1970",-0.00151193683336825,-0.010509701675576,0.00529083661088747,0.00144517657820198,0.00226521694457471,-0.00331993766272087,-0.00739836932507931,-0.00638510573678353,-0.0143098562965259,0.0116697308327325
"1971",0.00641058578261045,0.00600318488553353,0.00789471558180299,0.00937943324935464,0.000837096658570013,0.00104693562310043,0.00853763510978589,0.00975766032359582,-0.0104802161161337,-0.00842948025412049
"1972",0.0114352864229668,0.0119351284571998,0.0496083980105246,0.00428879967766527,-0.00259312017041191,-0.00161617369181166,0.00752501218603974,0.0254535415487167,-0.0219636943838234,-0.00134235562090357
"1973",0.000545564083670236,-0.0131553260493088,0.0066334938403172,-0.00830366106145441,0.000000222181523179543,-0.000371689025722599,0.00773539318186689,-0.000919212938876091,-0.00452691267435068,-0.00896049769793583
"1974",-0.00346932209294692,-0.0022981338042718,-0.0263591222859495,0.000956769778817756,0.00311008661194134,-0.0000952802618869875,0.00119104439273232,-0.00897167498105034,0.000624155138222893,-0.0144666273901938
"1975",0.00631646646654982,0.00691093261422671,-0.00507616704416425,-0.00884279962471601,-0.00142433232135286,0.000285772201556789,0,-0.00789205999746312,-0.0216538939435582,0.0027524450020886
"1976",0.00400285575852322,-0.00388928135408584,-0.0127551766473719,-0.0122983401599205,-0.00646180359025295,-0.00305277302064422,-0.00422989986863631,-0.0138047356795331,0.000819710348668234,0.000914806340723828
"1977",0.000935263196630842,0.000229571209025003,-0.00344507833317453,0.00634767027416094,0.0114874557073363,0.0064112771019198,-0.000796695999289776,-0.00450740184159026,0.0281216243571611,0.00457041564431049
"1978",0.00314734228992331,0.00459258558472952,0.0077785257997729,0.00266869957139138,-0.00918574538647354,-0.00408837855077049,0.00451712556574346,0.00762622770692656,-0.0222183055482137,-0.00955414996961046
"1979",0.000980544498284663,0.00731413551588167,0.00600353515840601,-0.000967760433172704,0.000674193791925459,0.000095089872978571,-0.00251287600433892,0.00614935041139897,0.0143038386230658,0.0050528032285897
"1980",-0.00107731966699109,-0.0115724258969453,-0.00511502075947623,-0.00193772742416842,-0.000842547083976131,-0.000381686645765655,-0.00517112507250328,-0.00376107748513255,-0.00481971612977761,-0.00319922509623971
"1981",0.00112757315679235,0.00367301943404708,0.00856894304637112,-0.00266923656472817,0.00236054191206425,0.00162378921036677,0.00399861295068238,0.00283145744469482,0.00152464573991029,-0.0183402430648723
"1982",0.000244928081769569,-0.00091496170809513,0,0.00827242849494958,0.00487762865034891,0.00209756713614784,-0.00610634108977437,0.007058770137363,0.0250739057056308,0.0107426411771041
"1983",0.000636467504940397,0.00228929706553838,-0.0161426778798385,-0.010617825442453,-0.00251047790809267,-0.00114162844342258,0.00373955022001637,-0.00420568471098648,-0.00366906609881124,-0.00415900323180507
"1984",0.00577379399873368,0.0139333666414849,0.0138170078239683,0.00536603983922079,0.00276836019943927,0.00114293324852799,0.00479068311232211,0.00375408243366948,0.00876808394297024,-0.00510438663375412
"1985",-0.00160546075136148,0.000225466850489298,-0.00596262356279809,-0.000485019295579647,-0.00635864402590869,-0.0026642243195012,-0.00622468384319896,-0.0021035855032594,-0.0119078919102679,-0.00513052706809547
"1986",0.00175424303083771,-0.00427935381304312,-0.0102828965630679,-0.00169915291614597,0.00522072896543424,0.00181258797243689,0.0027985169066651,-0.00960406461843266,0.0103800228712174,0.00843884767950143
"1987",0.00535068181130449,0.00814304049672132,0.00779218677140614,0.0318503043822655,0.00603098685827885,0.00200029542635161,0.0073091489128303,0.00946044937102108,0.00461429562411375,0.0106925542322909
"1988",0.00280623193532947,0.00830132168516373,0.00171818221583875,-0.00824702731171767,0.000832649059381074,0.00114016700776221,0.00290242219657078,0.00164013031043941,-0.00242653611601129,-0.00873962635098224
"1989",-0.000723895020825593,0.00356062305733085,0.00257322994860032,-0.00641479020658531,0.00831962067969183,0.00246834807360785,0.00276217792037192,0.00233920669682197,0.00234554771657081,-0.00464030806755011
"1990",0.00255918126719967,0.00421262020531654,-0.00256662543117403,0.0126731486018372,0.0027226012483339,0.00170409117539139,0.00747764114394878,0.00210056463584052,-0.00190668231686641,-0.00233111440108369
"1991",-0.0021187410871929,-0.00684483670413549,-0.00343037594504048,-0.0200707596805669,0.00789917095677062,0.00387594385062728,0.00286437102419268,0.000465675427002932,-0.0264849157177869,-0.0457943004701402
"1992",-0.00695001404496731,-0.00111152699211581,0.00516351249071656,-0.017108352772581,-0.00583405983455498,-0.00245220517123335,-0.00363546916871216,-0.000232681506243004,0.039871563287204,0.0205680919931677
"1993",0.00646362803478517,0.000222468979377055,0.00856160675515216,-0.000245136064642826,-0.00971211135717376,-0.00444445001487215,0.00351862867990138,0.00651899056959704,-0.0123520584602493,-0.0211132512505544
"1994",0.00386318956561404,-0.0017798272112558,-0.000848881120165457,0.00269749365191507,0.00390674675084712,0.000379925282137039,-0.000909449312037625,-0.000231006467610761,0.0103352701957204,-0.00588237341865872
"1995",-0.00110625744319925,-0.00401268247262065,-0.00254871356243547,0.00171175574720861,0.00836136093617945,0.00351311167125301,0.00156016347367749,-0.0115689350087295,-0.00386834859677898,-0.00295853949162506
"1996",0.00163711544125911,0.00492373035329186,0.000851585915721875,-0.00195322788918806,-0.00582934765593812,-0.00558247505900389,-0.00519074966313493,-0.00304316798334092,-0.012512918860362,-0.00247276535029672
"1997",-0.00668268171915154,-0.00757230180445279,-0.0161702493860182,-0.0146769573009685,0.0122224104596051,0.00333014604106219,0.00443515495899338,-0.0150271645268342,0.01179759678406,-0.0173525206683872
"1998",-0.00067754159772504,-0.00875208273382988,0.00519043226442739,-0.00943362312775897,0.00514013969391236,0.00369823682057935,0.00337683840101577,-0.00142999598049365,0.0208153655278578,0.0070634753146015
"1999",-0.0160311027644319,-0.0115464113696251,-0.0154905138125769,-0.0147873760253405,0.00730500682423241,0.00453540358024362,-0.00233010800585787,-0.0057291889447566,-0.00194604447168056,-0.0155310053935875
"2000",0.00506968271509689,-0.00366460694992643,0.00262216194503107,-0.00839478124684057,0.00410952563357037,-0.00169303460715986,0.000908252452273439,0.00432161015244703,-0.00228888608247602,-0.00916028487234122
"2001",-0.0161614885797693,-0.0236780992112728,-0.00959018375992249,-0.0164187800287268,0.0135624334769908,0.00819662110598052,-0.00907341250293858,-0.00812815951179824,-0.00237911458273243,-0.00821792272696698
"2002",-0.00686927213053357,-0.0174241982691428,-0.0193660192966347,-0.0143452625404827,-0.00205862873769247,-0.00364416778694776,-0.0117723575543273,-0.0110869961852751,-0.0257218711959162,-0.0160538006646467
"2003",-0.00801975650262055,0.0119818465686925,0.000897649807543033,-0.00158769963061267,0.0123768159469626,0.00506450852575413,-0.00463278537708089,0.000974840123615373,0.00489551538504673,-0.00578939496770725
"2004",0.0196050739716911,0.0108927374970922,0.016780980490267,0.0229869720571783,-0.00901234210030266,-0.00690566244551638,0.022340582571762,0.00998316387807985,-0.00591561563938092,0.00582310723543245
"2005",0.0247287344996472,0.0210822788000355,0.0159715707239061,0.0136662620944838,-0.0177933798526679,-0.00563815664907474,0.00897492512957521,0.00867884129364382,0.00770110285379633,-0.00315774346202635
"2006",0.00425477247300798,-0.00145482026281596,0.00524013940097912,0.00700032384386806,0.0134457035683249,0.00368562223154156,0.00206280944766468,0.00320398783677045,-0.00330008678592986,0.014783378020544
"2007",0.00459990178611669,0.0043939026707851,-0.00260645922823621,0.0139031172125148,0.00135073400046459,0,0.0164669365828638,0.00816533964232069,-0.0193429821210155,-0.0182101106723288
"2008",0.0013497201397632,-0.00368400542066438,0.00174217247224173,-0.00914177119335313,-0.0198348662617323,-0.00828539003073636,-0.00506238967346717,-0.00119109410964247,0.0016880941353683,0.0100688091195851
"2009",0.0000961054470451916,0.00670218787615751,-0.00173914258590324,0.00230675197375674,0.00544276493884444,0.000722448084400362,-0.00411287299241825,0.00166963050524305,0.000266090123578033,-0.0131163498056155
"2010",0.00322462402471646,0.00114777044022385,0.00696861846991825,0.00792612556565708,0.00371122344310493,0.00133051478969315,0.00387194590717344,0.00428555985254087,0.0182673144879129,-0.00106324961847593
"2011",0.00134343386608782,-0.00802569121672625,-0.0103807193670878,-0.00608815914227478,0.00747513173544689,0.00341556411750288,0.00437095830723577,-0.003793274039531,-0.010101924408222,-0.00957959621759008
"2012",-0.00536588770145519,-0.00970869484683445,-0.0122376104636792,0.00204180771917417,0.00271267326642288,0.00113487027341463,-0.00102411285322268,-0.00309362514193323,0.0134600072747426,-0.00107467628639846
"2013",-0.00992284128898646,-0.00723641500154037,-0.005309771497926,0.000764121294750231,0.00190973468909461,0.0011334052212022,-0.015376573774756,-0.00763887327641077,-0.0140624569634321,-0.00753093793412274
"2014",-0.000535398755257765,-0.00493761491896405,0.0017795664081548,-0.0132348375507283,0.0111180217061335,0.00509507395214337,0.0123631975872294,-0.00192472927651,0.00440218340549059,-0.0119242345282613
"2015",-0.0180596520025051,-0.0300094287272753,-0.0115455050279215,-0.0177972581442536,0.015709013816132,0.00610118069361443,0.00334255766406311,-0.0060256084099366,0.0150771473513824,-0.014262180473698
"2016",-0.00941905009371058,-0.0107186118468209,-0.016172448230189,-0.0042018427693199,0.0180168818106923,0.00671791665909605,0.00730289367836234,-0.0033946369316924,0.01139896343526,-0.00946031160562877
"2017",0.0124613259478481,0.00935732841357972,0.0146116991680718,0.0216247652608099,-0.00197496927268881,-0.000185343497561719,0.0129737000384147,0.0167884993814513,-0.00589141890646971,-0.00617957602536812
"2018",0.0177449915337795,0.0153693915787678,0.0126013006670609,0.0170364858573335,-0.0132427935495468,-0.00407858087117219,0.00565027481732594,0.0107678669166,-0.00420852014085715,0.00395698354185292
"2019",-0.00801348921540423,-0.00624664794509755,-0.0106665964435301,-0.0032995502253671,0.0109523357482115,0.00493272448519821,0.000374884061584257,-0.000236501563094849,0.0113851990445886,-0.0016891660869599
"2020",-0.00783370897206803,0,-0.00359401380102675,-0.00814868548114678,0.00572236823314443,0.00351965614828553,0.00549184645125034,0.000946841463282722,0.0110864401997877,-0.0219966048061198
"2021",-0.00281269552093732,0.00435170824873365,0.00811548951632735,0.00872911991823933,0,0.000923125304537198,-0.00260698336835075,0.00828042562192088,-0.00337376861291772,-0.00403703159616031
"2022",-0.00603724168070185,-0.00192568428079432,-0.00178872584237433,-0.00559937306810809,0.00758586814819395,0.00461021084760271,0.00659620557142304,0.00375401650079854,-0.00160801450209835,0.0110017664138224
"2023",-0.00916039811582126,0.00603006822401086,0.00716833668762784,0.0023035981737054,0.015735252679467,0.00853567863631177,0.00135974860527299,0.00186990886703842,0.0251759004392991,-0.0137458120305932
"2024",0.0131142123743626,0.0141451506021539,0.00889668925126719,0.0084268554257465,-0.0127487839976435,-0.00737115180670289,0.00851983311953108,0.0177322472143784,0.0130642878606864,0.0191638030508074
"2025",0.00213256165105324,0.00732860151693537,0.00793676921390629,-0.00151942726812648,0.0132892135161327,0.0022918799200895,-0.0078352298054658,-0.00802396531516991,0.0137120473484831,-0.0136752043521947
"2026",0.00504800370438074,0.00774454021818838,0.0017496976220186,0.0220647226386592,-0.0115588162154665,-0.00475654000088566,-0.00148101570764336,0.00762652963222243,0.000241594208734153,0.00635480048784021
"2027",0.0148709698501424,0.00302746061843395,0.00436675896542638,0.0191064458439032,-0.0035982257117213,-0.00248177666628857,0.0195255615229522,0.00366951344949062,0.00804958525196198,-0.00114808995632198
"2028",-0.00548291477207985,-0.00510777636618742,-0.00347819011201866,-0.00754800265325783,0.0139181457385533,0.00654179813873301,-0.00206079433530293,-0.000228162536320298,-0.00798530684376009,-0.00632181185090264
"2029",0.00234188305532745,0.0151689577891714,0.011343537195549,0.000490602953983288,-0.00304232390759085,-0.00228847712849944,0.00983842117250422,0.00617161005327116,-0.00998152596035917,-0.0034702855386991
"2030",-0.0131905339336503,0.00137955778866994,0.00172573225129136,-0.00539467579052755,0.00156312729825392,0.00137648065931151,-0.00132278672002706,-0.00477082861059774,0.0114643794042504,0.00522343606937192
"2031",-0.0128244762826306,-0.0197427892002255,-0.00172275923012666,-0.010848177406077,0.016348523594903,0.00769665657609253,-0.00710595185529461,-0.00890204677591611,-0.00787784553251047,-0.0144341619889924
"2032",0.0092437060515671,0.0170957496702793,0.00862828396990811,0,-0.00658023801100815,-0.00354636002143349,0.00169843986390683,0.00967304162213156,-0.0215523905615361,-0.00468652079010523
"2033",-0.0125749521160368,-0.0161178298300321,-0.0171086899203288,-0.0274178354577719,0.0177370174688136,0.00875991477482585,-0.016348009361679,-0.0177918771427142,0.0222755461696662,0.0241318147701892
"2034",0.0123840801891102,0.0109992911447581,0.0104438667760076,0.0179394599334275,-0.00377609267078305,-0.00125029896091466,-0.00320059474134904,0.018810755026329,-0.00834345099255041,0.0137930332837239
"2035",0.0144611365900045,0.0217591377897821,-0.00172275923012666,0.0188823678426122,-0.0211656615113055,-0.00843673428352854,0.0092623974511814,0.00866215733932818,-0.0111909412055373,0.027777866916868
"2036",-0.00380780770882272,-0.0124601084456105,0.00517710243223668,-0.00494201883415069,0.00170882685908968,0.00164691945992534,-0.0029368277333417,-0.00949172499509388,0.00437834768166012,-0.0220628612013305
"2037",0.0100951526763737,0.0137644898186378,0.00858368031480805,0.00595976468879389,-0.0109792450834173,-0.00365364574232219,0.010431904733188,0.0182520306259593,0.00172724951920977,0.0135363096736323
"2038",-0.00276534935693695,-0.0153882017800211,-0.00851062780643919,-0.0170327147414101,-0.0177017226978684,-0.0111847890216122,-0.0263571768651385,-0.0100825445916307,-0.0258642086717776,0.00278243448269144
"2039",-0.00447594336865653,-0.00390695323083101,-0.00944206711345663,-0.00150683510925509,-0.0016036735729722,-0.00046313815666188,-0.00474048442162922,-0.0140336162060201,0.00446728763037174,0.00998887909743806
"2040",0.0106531413146242,0.00946004322333671,0.0129982034637515,-0.002515191243597,-0.00795399578550104,-0.00250460335208236,0.00350942776571816,0.00367325744661295,-0.00587393649196843,-0.0126373600584188
"2041",0.000580509537600138,-0.00617149274079309,0.00171089938433133,-0.00731214048748963,0.001850355300137,-0.00037164598429984,-0.00212289485421602,-0.00251615515651882,-0.011817346063836,-0.00779065618397379
"2042",0.00961672535010027,0.0200091043333213,0.00683165210234637,0.0213361330835264,-0.00330875459258806,0.00037178415638861,0.0107645477976359,0.00986018884986617,0.00230627829503716,0.015142982519029
"2043",0.00411645878802513,0.00338229312390137,0.0118745774357853,0.0114398052731011,-0.0102686798208361,-0.00334776670766868,-0.00544899981915692,0.00681193957708115,0.00545429539643072,0.0110495723323076
"2044",0.00157325253626195,0.00247197679955757,-0.00083833192129934,-0.00221283418380602,-0.0150559976112664,-0.00709081454603699,-0.00286387750642525,-0.00270602778408391,-0.0166977534319948,0.000546553163430996
"2045",0.000094946054344458,0.00403488063885282,0.0176174487796397,-0.000246292541873694,0.005940173904041,0.0047922270352927,0.00849166971079884,0.00248745837256559,0.00284453059487055,-0.0120152404922721
"2046",-0.000713503370640467,-0.00178605919309172,0.00741986502736891,-0.00419038919676973,-0.00661348883746193,-0.00252482192267622,-0.0190688921430249,-0.00383477367904017,-0.00343814692928124,-0.00331676100198663
"2047",0.00600027819110571,0.0134198692748879,0.00900153073077781,0.0066830349572895,0.00293243497081908,-0.00056262011773478,0.00921494646446841,0.00543445229120332,-0.00569262539774673,-0.00388247916964912
"2048",-0.000141980494039906,-0.00441404513601862,-0.0056771720541543,-0.0100810148175671,0.0114584239441351,0.00459691302882614,0.00787959030501639,-0.00180156025034539,0.00130118842211302,-0.00668153796059567
"2049",0.00284086636192948,0.00620692671330225,0.00489384199722331,0.0144062202854209,0.0131260978445302,0.00662959819529929,-0.0188629838315296,0.0051894623034745,-0.00147273672355541,0.000560530484758237
"2050",-0.000849764754779603,0.000660851057200817,-0.00243518193699088,-0.00195873323608975,0.00431866387483337,0.000927811475744944,0.00215010379218339,0.00246903314169078,0.00381741273959024,0.0151261328873129
"2051",-0.00118130576317454,-0.00462344272482473,0.00895061935669061,0.000245398068674074,-0.0136680679555031,-0.00593119882220861,-0.00845670148555244,-0.0033586401096698,0.00319795168188297,-0.00827820277748603
"2052",-0.00340629639497414,0.00176967362363434,-0.00403229699012431,-0.000735792862886497,0.00840772188679995,0.00354263726902926,0.00712881305244673,-0.00292071219445356,0.000775428620660046,0.0111296806566363
"2053",0.00631357661855581,0.00154544189349326,0.00242893434596714,-0.00147291780585745,-0.0186263626151315,-0.0074440857533361,0.00391793310710953,0.00856236894259044,-0.00413226569792469,-0.0143092756386252
"2054",-0.00410406519539941,-0.00859793104031126,-0.00484640689799709,-0.00762055888744018,-0.0036256353572659,-0.00215631204077593,-0.00264373077451852,-0.00513854076202436,-0.0018153440525589,0.00614179367706202
"2055",-0.00421578792017685,-0.00378010976708776,-0.00487000894293144,-0.0108990134777653,0.000316117657937598,0.000751526885606424,-0.00833166724013623,-0.00763525463859704,-0.00311769288024866,-0.00887895921922588
"2056",0.00109419579407111,0.00334821422748166,0.00570958635826835,-0.00150257146017962,-0.00126481906092957,0.00056365638226441,0.00330998451742026,-0.00045271488234444,-0.000955616358651601,-0.00391931914536592
"2057",-0.0140644860916124,-0.0180202091429446,-0.00162207132352732,-0.0152997942376961,-0.0220919210041354,-0.0102272405190421,-0.0304491060042471,-0.0185646404204682,-0.0273043391304348,-0.0123666170244006
"2058",0.00414463457385894,0.00385148148507097,-0.00324932462255556,-0.0038205205176266,0.00923056352603258,0.00464516605786636,0.00889799186866913,-0.0129179130731153,0.000983372063442012,-0.00284572097699964
"2059",-0.0162220466894625,-0.0243735899007139,-0.0146699835596452,-0.0222451358907576,0.0131578799392726,0.00424628872062516,-0.00492843704728796,-0.0170600733274772,-0.0049120567570593,-0.0131278504276504
"2060",-0.00234176890479965,0.000693870555953824,0.00909843539001631,0.00758378599620735,0.00728542818162814,0.00178498456262077,0.00143371882243803,0.0028528779783028,-0.00601326523089696,0.00520530925471774
"2061",0.0127139373751517,0.00809062406724048,0.0221312457214757,0.00622890468572401,-0.000707731938503153,0.000937533872415353,0.016529909917113,0.0109058883929571,-0.000270871331828459,-0.00460298819676297
"2062",-0.00613196685625439,-0.00710853827792268,0.000801765756319961,-0.0121229003937716,-0.00306801824997527,-0.00149886106752262,-0.00371325325852867,-0.00257988494799288,0.00144505056498345,-0.0202311155214705
"2063",0.0133603523328292,0.0145495361240835,0.00400644936891292,0.0120105086627447,0.00962765514343555,0.00347170546057396,0.010924190906092,0.00940527028600946,-0.000631304129634969,-0.00118004618052503
"2064",-0.00297241557623917,-0.00409723169282117,0.00239436867938236,0.011609704665535,0.00828482382528439,0.00205781720534204,-0.000890099460170823,-0.00652231946013015,-0.00541466483917807,-0.00708803408364778
"2065",0.0120215261647645,0.023771352202008,0.0159236110905605,0.0244836406363576,0.0193026756186563,0.0114793325963838,0.0197227681509606,0.0192260062619907,0.0195989839361128,0.0273645963994336
"2066",-0.00456142145579663,-0.0136190829727528,-0.0117556625939653,-0.0169280188439819,-0.00509577854296051,-0.00470569843346558,-0.00149741793333891,-0.00253031379261115,-0.000711951569494884,-0.0167920756911898
"2067",0.0088270454358037,0.0251245767472523,0.0158604960865336,0.0149406407584391,0.00527447408338211,0.00407875070148189,0.0242440354084161,0.0197232849749041,0.0113990470086467,0.0135453445761553
"2068",-0.00194866696371443,0.00507830446234947,0.00468370259880579,0.00299400819472151,-0.00121654327272447,0.00129281069031384,-0.00146416625784362,0.00136204239417292,0.00633971119133592,0.0116211714476675
"2069",-0.0056189538469571,-0.00175759599771141,-0.00233092328065021,0.0039801411275513,0.00966890025919342,0.00304303257071825,-0.00806471499463135,0.00702768289257572,0.00244989935733742,-0.00804142308010869
"2070",-0.0146539442751936,-0.00528145444245931,-0.00233639046276424,-0.0158575332361894,-0.00844540258079141,-0.00432102503957832,-0.0165174263863541,-0.00562815510085257,0.00139655232608882,0.00289521423429195
"2071",-0.00238144381096861,-0.00973456784936022,-0.0101485734425625,-0.0093151447637817,-0.0155892712664286,-0.0056317385065412,-0.00568228398753523,-0.00950858103682839,0.00653708690306587,0.0121247840176284
"2072",0.00228963198278098,0.00178725612513242,0.00394332148902876,0.00279547497246635,0.0124373864730987,0.00389969816730606,0.00342859369699822,0.00571446962333177,-0.00363703662182968,-0.0199657933908359
"2073",0.0121998090909283,0.00356834359857916,0.00392785425034448,0.0192601208409866,-0.00495999060904273,-0.0000929335745997184,0.0112645736668284,-0.00454552615656068,-0.011385346973498,0.0052385780379427
"2074",-0.00873948395201818,-0.0162222802500465,-0.0195618340941202,-0.00223781570973869,0.00214746810449329,0.00259017968321795,-0.00725901054707323,-0.0109588735374352,-0.000791173626373598,-0.011580737745951
"2075",-0.00353623637109524,0.00880951957286435,0.00399046178580975,0.0124596138096034,0.0131343443352374,0.00475911333512502,-0.000126548848109254,0.00738689869111675,0.0170683963727469,0.0181605695309341
"2076",0.00359739150110183,0.00806083185697437,0.00874404463177036,0.015013467263804,-0.0105953210432386,-0.0028510633113048,0.00668308347160584,0.00801998134326731,-0.00276815748733827,-0.00517835431905656
"2077",0.00673318488114472,0.00932914676635543,0.0118202730806536,0.0128517988628793,-0.00558372566438903,0.00129144514948831,0.0100200731367606,0.00727451515979238,0.0122311156508599,0.0127241223596799
"2078",-0.00264621510729601,-0.00154034061983443,0.00467292991916279,-0.00502764598010641,0.00838424096833434,0.000828914557561955,-0.0162452495894511,0.00157982217772856,-0.0049704429690558,0.00513984965216796
"2079",0.00337702341210533,0.00110187810271922,0.00155025010266652,0.020933522949617,0.000305453205501571,-0.000920558960303963,0.00277343120023099,0.00968854316538326,-0.00551201442156568,-0.0193180940344471
"2080",0.00442353003759166,0,0,0.00989859173509955,-0.012964406731139,-0.0040537327303577,-0.0175992245885058,0.00290137877355301,-0.00692823238132634,0
"2081",0.00545701148203626,0.00330269067815681,0.00154808323033562,0.000700312779423173,0.00146781083992198,-0.000276881819722297,-0.000639702825793731,-0.000445093174625488,0.0113369061016291,0.0104287728250716
"2082",-0.00452295046944451,-0.00548600563437585,-0.00695508923069765,-0.00583048283541698,0.00138887326706461,0.00203543917850535,-0.00281700050396017,-0.0131342568854391,-0.0071570405522372,-0.00458721091733771
"2083",0.00191298664087958,0.00882627107345035,0.00700380129364908,0.00445706037881233,0.00708782279096387,0.00295493050113249,0.00205446249379992,0.0090233782975182,-0.00607952932151745,0.00460835039256935
"2084",0.00448718411104121,0.00503046513697347,0.00463690215643719,0.00700601116824795,-0.000841221043894058,0.00055240628857911,-0.00589404937398308,0.00268258153532042,0.00865080376353022,0.0200688264583102
"2085",-0.000285328319723055,0.0017408684843716,0.00230746645775026,0.00788505904728987,-0.00497710425988451,0.000736090942920375,0.00412430905952799,0.0031213908324188,-0.00346531231049119,0.0106800103349713
"2086",-0.01150331784404,-0.0134692681474705,-0.00767450491202459,-0.0174873668515565,0.011464949481174,0.0020225703521799,-0.00526283974680231,-0.0115579666313371,0.00495522042037044,-0.00222466379608099
"2087",0.00913682154295659,0.0011009073722108,0.00309368710789393,-0.000936705578791996,-0.00882462740493306,-0.00183500462115227,0.00129039684475574,-0.000674756786301689,-0.00761243092755071,-0.00445924791956631
"2088",-0.0011913794132834,0.00769908530089825,0.0154200122003769,0.00586015596002931,-0.00452810226546696,-0.00211472436665627,0.000773517182882211,-0.00224998694542666,0.0057531031576612,-0.00727885080943291
"2089",0.00491422637328709,0,0.00759308914464207,0.0107202747777719,-0.0152661369812971,-0.0058034377388495,0.00296163656186899,0.00270629891828955,-0.0134338277023877,0.00338416449252255
"2090",0.00251633928038864,0.00545739215306695,-0.000753430339523353,0.00737842332054561,0.00430646084256225,0.0030575826721162,0.00179779769155908,0.00202442107324918,0.00729159259788115,0.01236644346353
"2091",0.0023206273259484,0.00434206937151016,0.00377069288524789,0.0036619973674894,0.00623701316752623,0.00351042670704049,0.00166608603414264,0.00606038540704579,-0.0140415222731023,-0.000555353763433186
"2092",-0.00415794175283313,0.00713370963992532,-0.0022540318886326,0.00387694678492845,0,-0.0015647289898334,-0.00268692679134586,0.00178504864305151,0.0201680578460488,0
"2093",0.00317871116290225,0.000429194712915359,0.00301198701189409,0.00158998412980105,-0.0137909703475212,-0.00461024486432049,-0.00025676470304048,0.00289523006805692,0.0086707706811624,0.00166675834314023
"2094",-0.00411454367611164,-0.00836734880661771,-0.00900884708485639,-0.0124743732133707,-0.0122557753188504,-0.00370491932281547,-0.0196354361319149,-0.00644010923906957,-0.00704891245510331,0.00665542577805445
"2095",-0.010020510195309,-0.00302889432991749,-0.0257577331730598,-0.015158302459654,0.00174963152417829,-0.000279244137630141,-0.0116507929893569,-0.00916407744585057,-0.0176608169394716,0.00771362090786609
"2096",0.0108415472823959,0.00802946493416057,0.0124418739327661,0.00606322365553336,-0.0134614432380247,-0.0054668729328935,0.00529771610610541,0.00248123967549962,-0.00343702297138437,-0.0010934787598561
"2097",0.00284740974939268,-0.00172225528584913,0.00460817972471861,0.00579513576567292,-0.00943557050011834,-0.00206034647418529,0.00263530917411336,0.00607538822656006,0.0090201271839383,-0.000547337882276788
"2098",-0.0114519210750519,-0.014880331184622,-0.0191130015585654,-0.0108321015573781,-0.00138376913506755,-0.00168892519429364,-0.0219449960472254,-0.0136432418663226,0.00280455745494401,0.00821473346996493
"2099",-0.00411687593032861,0.00678643904482135,-0.000779524420873701,-0.0123483283604426,-0.0171206800770177,-0.00488829848662264,-0.00268666785721372,-0.00680252310069007,-0.000524357638950534,0
"2100",0.00398955138283541,-0.00413154787440484,0.00156000929038846,-0.00141547941819009,0.0134373575814672,0.00425062409575849,0.0132022317088234,-0.00639280760151051,-0.00821968338387813,-0.0157523714176044
"2101",0.0131660918279448,0.0248909308995791,0.0233644367477643,0.0127568410812116,0.00270111467679635,0.00385657314625187,0.0152902370923467,0.0238971037725901,0.00484925947538795,0.00551868825165203
"2102",-0.00477266797699161,-0.00447382653370043,-0.0159817126514713,-0.00956378198702934,-0.0243247224145219,-0.00983846370306662,-0.0145364987796193,-0.0089764691612737,-0.00386068260190675,-0.00439071958871129
"2103",-0.00299131527106711,-0.00385183061309324,0,-0.00329733181367797,0.00259323716598736,0.000756946197094654,0.00292356157482709,-0.00181172689154518,0.00854400606486383,0.01047394718828
"2104",0.000190624758196423,0.00644468324428549,0.00618722625922885,0.00189052548368562,-0.00801058541000843,-0.00132371661034292,-0.00834739782156113,0.0111159353438959,0.0179039563318777,0.00109120500779669
"2105",0.0104276898438675,0.0164354009047265,0.00538044050122011,0.00990559505307886,0.00269168450091906,0.00340871615921068,0.0181719860050924,0.00964760835929424,0.00540537952624498,0.00599463697079994
"2106",0.00108373758736446,-0.00146992321994444,0.00458710449441968,0.00770678829372251,0.0200509892167593,0.00717195578900753,0.00826779623345253,0.00866672270801772,0.00298684929168802,-0.000541704379498187
"2107",0.00310674336494254,-0.00546799076422733,0.00837139211163618,-0.0101972435640756,-0.0167780554518283,-0.00674620195973985,-0.00299362770457967,-0.00837152798170682,-0.0000851016768919077,-0.00271010147902528
"2108",-0.000328514345499409,-0.0033832772081781,0.000754876993600551,0.00163917384500434,-0.00886661360086305,-0.00443375043921934,-0.00130545353181044,-0.000889042309883292,-0.0138699629136307,-0.0211955866319149
"2109",-0.000704329646047941,0.00297038630421809,0,-0.000701327141712893,0.00168795467547844,0.0021791371919293,-0.00209157082534084,-0.000444465104326053,0.00163951161998011,-0.00222107217221601
"2110",0.00291245192524792,0.00571195251883672,0.00377069288524789,-0.0035087546648277,0.0139860940918837,0.00595658766641538,-0.00458480889179014,0.000222466911058872,-0.00335975183735771,0.0122427460883201
"2111",-0.00238854025142221,-0.00946561471426122,-0.0022540318886326,0.0032863106565002,0.000415127333581289,-0.00225534209933964,0.000263032407725738,-0.00556091757759891,-0.000777975611064519,-0.010995183959485
"2112",-0.010751866567927,-0.0205990265379452,-0.0128012432045435,-0.0159101191492924,0.0171098036902044,0.00621695995093963,-0.00605157483764229,-0.0138667516494407,-0.014619325512445,-0.0194552740661222
"2113",0.00949217900381671,0.0125760487271396,0.00686513081030315,0.00023770628200892,0.00228647294068063,-0.000561732280637939,0.00754465374270619,0.00249474600815924,-0.000175621098213563,-0.0136053739085655
"2114",-0.00112824744433726,0.000642213034935057,-0.00227291897580095,-0.0130735460327484,-0.00244421505826697,0.000936615553712272,-0.000656826724706905,-0.00610849910592204,0.00114143472773232,0.00517234311863457
"2115",-0.00621289716948115,-0.0113415748924282,-0.00911145380557776,-0.00963373012513336,0.00220524189005067,0.000561687534633037,-0.0107797891596851,-0.010243609128223,0.000701640081607779,0.0125786219037087
"2116",0.00203663680976174,-0.00692650084535951,0.00459758647233666,-0.0038911736324827,-0.0107477209577789,-0.0044125712690477,0.00970135712434206,0.00184018619519399,-0.000876406676185937,-0.00225858023963132
"2117",-0.000992822855492959,0.00762850307570617,-0.00228827270453691,0.00390637401203686,-0.0139517087347096,-0.00696262712096585,-0.00816023258615473,-0.00114795332423157,0.00403507894736843,0.0118846210882944
"2118",0.00264965084275826,0.00865243332069277,0.00382266717333835,-0.00510701151507509,-0.0160751647511868,-0.00852744126205229,-0.0120751512916616,-0.00459693495765356,-0.00716407484854154,-0.0128636462591393
"2119",-0.00844675409231832,-0.0113660975154501,-0.00685444403629143,-0.0151553200748639,0.0130189960110318,0.00487348478994054,-0.000940590572775069,-0.0092356097231443,-0.00703980118831227,-0.00906514926579005
"2120",-0.00171319448303697,-0.0140997674892698,-0.00613517916579243,-0.00446754918736336,-0.0121795674500408,-0.00722774380306523,-0.0120997231167856,-0.014681760823089,-0.0053172458460562,0.00457409782496465
"2121",-0.006149501635203,-0.000439960035613307,-0.0054011990311793,-0.000249374866120977,-0.00110541817455689,0.00143713876854723,-0.00204130885153586,-0.00402115269649617,0.00294014616785709,0.000569144195399662
"2122",-0.00014403864244561,-0.00506268067358207,-0.0100851223396964,-0.00598483460768207,-0.00791697127135904,-0.00325222831513927,-0.0072276963879494,0.00522474112848736,0.00222084036599446,0.015927265450697
"2123",0.0119934055258697,0.0250001001972269,0.0164575892232284,0.0145509002263613,-0.00875243531061343,-0.00383877086143203,0.00714275223633409,0.0181905243223563,0.00850912072327614,0.0039193191453657
"2124",0.00322347989562166,0.00215809196698791,0.00462586037416601,-0.00494565713090578,0.0210352524706827,0.00789963892676626,0.00791032739360853,0.0025519553436244,-0.00457019691132188,-0.00892358463847098
"2125",-0.0076549319033079,-0.00969178464949516,-0.00537218280263041,0,0,-0.000573924890084676,-0.00189417506442113,-0.00485990087500454,-0.000264868439610377,-0.010129466925154
"2126",-0.00428530613150435,-0.0108744027842839,0.00308661032363911,-0.0111830429948711,0.00161093331226692,0.00239138681610096,-0.00515188603499095,-0.000697477704375227,0.00441579075114928,-0.00454797665417239
"2127",0.0054516111746894,0.000659646066439201,-0.00461550053206694,0.000251408685866261,0.00787186227892223,0.00381602963410765,0.00844916739610913,0.00023249729984598,-0.00360505573889769,0.00285547202898218
"2128",0.0016170291002271,-0.00131842244070157,-0.0085006106411547,0.00603045477594177,-0.00772599013082187,0.000570706647145869,0.00621614502452572,-0.00302466040572447,0.00467700317684439,0.00284745874768899
"2129",0.0103995414550757,0.0127612325392066,0.000779268804176114,0.00924049775159075,-0.00490924203363374,-0.000760141330842679,0.0138330220772367,0.00560090261532276,0.0129117437489985,0
"2130",-0.00443921211986054,-0.00391050886127831,0.00077889615001081,-0.00866126325682326,0.012843110962758,0.00532408259158501,-0.00649121246336593,-0.00359054688420024,-0.00173427852930974,-0.00908585572589227
"2131",0.00512308228588298,0.0233370157318404,0.0155641824732395,0.0144782566832244,-0.0204063874059022,-0.00841634344670938,-0.00986647565659937,0.0101271261706755,-0.0128561845155615,0.00343846653051139
"2132",0.000707889105712622,-0.00149182817427473,0.0114942803151841,0.00984274858260092,-0.0060007980508624,-0.00305157024931146,-0.00484798903136252,0.00373081212335546,-0.00659978886483448,0.0119930413004823
"2133",-0.00726285654561276,-0.00787788916306964,-0.010606154653813,-0.00706648201913584,0.00862432424597892,0.00296557399867203,-0.00562475107829319,-0.00766574983207635,-0.00265748075699779,-0.00677197507159488
"2134",-0.00304060994019639,0,0.00200103132957596,-0.00343622302056601,-0.00350563509320168,-0.00247991010683646,-0.00947426990540701,0.000702457821972535,-0.00133221427594676,0.00113634815293406
"2135",-0.000190455219946428,0,0.00460813632443147,-0.00942705330958582,-0.0112407831536813,-0.00478052381328287,0.00485159893442111,0.000233706364646036,0.00106720026561358,0.00454040856141935
"2136",-0.020970264790056,-0.0335599003210861,-0.0252292730223584,-0.0222891232222857,0.0264689165826095,0.01162462445579,-0.0160021330837393,-0.0240877365798423,0.00453093469315813,-0.00451988643037415
"2137",0.00209318055407004,-0.0074896524076945,0.00470589133525623,0.0148566487028694,-0.0069329376941536,-0.002754075836507,-0.000420635146351822,0.00311530018104644,-0.00619082869019183,0.0215664003574805
"2138",0.00801550184790512,0.00548819318490334,0.00702570017775339,-0.00075716536810666,-0.0134978066494434,-0.00522650794587254,0.0152873253068826,0.00334426851179082,-0.00347067713435945,-0.0122220558958132
"2139",-0.000915647490750127,-0.000227653591741039,0,0.00479913652658115,0.00328621983791377,0.00354737282806661,0.00221046029086502,-0.00214286224346794,-0.00196464541977193,-0.00168738161556348
"2140",-0.00284571183764359,-0.0245676739128906,-0.00697668408712249,-0.0279034215580072,0.0185351453698013,0.0070695827125391,0.00454832904323244,-0.00978257546353978,0.00268428771144791,-0.0326760730635546
"2141",0.00628860621402971,-0.000932719458550557,0.00234185052997038,-0.0149986820313885,0.00939444148527824,0.00265636878244901,0.0153680285100168,0.00192770770260053,-0.0116008925861304,-0.00582415211058229
"2142",-0.0167772092911302,-0.0147060330683445,-0.0412772163279491,-0.0343921490548758,0.00863668035059884,0.00397387690431406,-0.00527036775888401,-0.0264551605399085,0.00297936072626648,-0.00468652079010523
"2143",0.00180891447092368,0.017531390672153,0.0121852497783699,0.0193038510465173,-0.0197026593331493,-0.00697395543830071,-0.0047545809418934,0.00963423243949735,0.00243050688380619,0.0117715903659563
"2144",0.0125913136607858,0.0419092284953779,0.0160513219808289,0.025339829434893,-0.0158580440142241,-0.00692768806597266,0.00696132250018788,0.0200635076594387,0.00116735810733348,0.00465380499809842
"2145",0.0110373200583094,0.000670441928616539,0.0134282140351618,0.00676402363434625,-0.00310192419726962,-0.00267615721485592,0.00149116219723844,0.011513506151168,-0.00448470722907357,0.000579150118952709
"2146",0.00433809417615416,0.00848590908404367,0.00623522067509064,0.00180884375547286,0.00328446582569453,0.00316212426405627,0.00270693198383531,0.0075886414664883,-0.00225245521673045,-0.00347241290050826
"2147",-0.000332200687430673,-0.00465010480117622,-0.000774549255890156,-0.0113490125856492,0.0105973516969335,0.00382052948366529,0.000945085681824498,-0.00282415821184878,-0.00523743914100483,-0.0116142449742631
"2148",0.00802427792832816,0.00912117231600473,0.00387595902478099,0.012522860485618,0.00690539324665296,-0.000380213090200865,0.00714761992018897,0.00991273794884528,-0.00363110008601675,-0.00470034876032666
"2149",0.000847921626159431,-0.00352730129228995,0.00231644940071662,-0.0012883280471031,0.00516435205546273,0.000095210025461423,-0.00388341154355909,0.000467476408399392,-0.0101129735766586,-0.0053127963211177
"2150",0.00051781680630647,0.00309737719400838,0,-0.00645006511597457,-0.00421167432095537,-0.0019989790145164,0.00174781257553458,-0.00186918828344673,-0.0271514491090392,-0.0160238240596492
"2151",-0.00395133256077373,-0.0037495559283961,-0.00308155193037907,0.000259817874078028,0.00541353912968945,0.00276579040138336,-0.00362323792843022,-0.00397831585359998,-0.00312198684357579,0.00422195857957752
"2152",-0.00179454427556747,-0.00730578106675084,-0.00463671042927738,-0.0142784448195653,0.00622625055415971,0.00123643005079099,0.00282835783119739,-0.00258432343014736,-0.00540950919399696,-0.0144144029424824
"2153",-0.00563012948085828,-0.00289908507749503,-0.000776501056808598,-0.00974450919134096,0.0124579098843891,0.00408506775448614,-0.00711799171043326,-0.0110722334831893,-0.0044847422380323,-0.00853139209343812
"2154",-0.0103719696462927,-0.0118541989272615,-0.00932388043902888,-0.014361677122981,0.00247730481016939,0.00094584914625373,0.000270408680357548,-0.00261999714165895,0.00977663165385545,-0.00799018329028789
"2155",-0.00581734547684576,-0.00792224497191951,-0.00392164364734526,-0.0188882648227411,0.0053549045701502,0.00330840583879377,0.00216364976784122,-0.0028659455205895,-0.00465113440248954,-0.0192069322486307
"2156",0.0122829505503039,0.0134611550974038,0.00472459010784543,0.0101759897054439,-0.007292665348688,-0.00282646253560215,0.0018891775953116,0.0124547492516616,0.0015258058218024,0.00821227311896955
"2157",0.00687929340964133,0.00225138335595965,0.00391839936936011,0.00980122496236402,-0.003714391664147,-0.0014168779735636,0.00511793584016984,0,0.0014283089343452,0.00313291822478545
"2158",0.000237081860148036,-0.000224557929096481,0.00156133982082007,-0.00997573800282281,0.00770489537259067,0.00113501480656431,-0.00375202802742691,-0.00260205383224554,-0.00855758312365851,-0.00374779901424127
"2159",-0.00151783958083596,0.00629068257995868,0.00779412651414724,0.010893097792551,0.00739960684470287,0.00585934021010881,0.00645615826978108,0.00308343118449916,0.00632974987042534,-0.013793109233514
"2160",-0.00337285758876904,0.000223076290120527,-0.00386696602215908,-0.0167024739254332,0.0105266496257099,0.00304814633611228,0.00494433283022055,-0.00425630330985316,-0.00791005432192893,-0.0165288315302095
"2161",-0.00195424274536748,-0.00267854462952677,-0.0015528543333122,0.00356167573403332,-0.00793199371555597,-0.00515921933871044,-0.00518596124720383,0.00403676162054611,0.00201729110503912,0.00581769849731795
"2162",0.00329537621659215,0.00671441039215237,0.00622082402913393,0.000272908917342551,-0.00750610562896792,-0.0038660613278666,-0.00427761750200728,0.00496717436646299,-0.00364296814577625,-0.00385605447913029
"2163",-0.00818780968077337,-0.00111153666694763,-0.00309114028618496,-0.00873347580982597,0.00887799448717219,0.00350245720206699,0,-0.00117694266281965,0.00442604637736932,-0.00064521886644664
"2164",-0.00191982918471967,-0.00400622973571596,0.0031007250623416,-0.00055072243045351,0.0131182747610914,0.00396196104849134,0.0034902171205089,-0.000942190366558626,0.00249068878715097,-0.0038734139922495
"2165",0.0125992460076547,0.0118436799525619,0.0146832420699354,0.0168044749183711,-0.0123854756636845,-0.00413429732060377,0.000134093398754809,0.00778260371318273,0.0102245482995786,0.0213869496870762
"2166",-0.00902325009125804,-0.0136927056314117,-0.0175171734578576,-0.0219454295145474,0.0158792722323575,0.00660450787451983,0.0066878327624178,-0.0142752679097928,0.00510784141971388,-0.0133249515791739
"2167",0.00119815221340636,-0.00582164161812793,-0.00620147120342451,-0.0155122246517335,-0.00545100687145139,-0.00037503707765818,0.0014618170418299,-0.00261192343189698,0.0140221905887035,-0.00321539024234307
"2168",-0.00124450789912522,-0.00292804652528778,0.00780012164942057,-0.00168833317446659,-0.00322359295521513,-0.00262505841880201,0.0019898949845325,0.00166641918655763,-0.0082598515081207,-0.00451613365891079
"2169",0.00364240330961119,0.00158117087591081,0,0.00140908769195658,0.00234472034173416,-0.00103437426638897,0.00569381876090547,0.00617849155918604,-0.0000936084587908059,-0.00648092618506435
"2170",0.00558664131750763,-0.00360844368376156,0.00232208093708408,-0.010976612862828,0.00451768543218112,0.00178815107276287,0.00750524729416746,-0.0002358114224561,0.00262048671259696,-0.00391384098282155
"2171",-0.00289660495953892,-0.00565873528825733,-0.00694983114135628,-0.0108140188744875,-0.00787013321736374,-0.00159702316106203,0.000783736487734554,-0.00519736207210519,-0.000186651736768018,-0.00523909389894606
"2172",-0.00790531197844702,-0.00956063419133557,-0.0108863997623718,-0.0123703548731541,0.00987505653173248,0.00611572807596805,-0.00548443389567332,-0.0047496176030023,0.0134441414112207,-0.0111914887418054
"2173",-0.0208814645735191,-0.0216042885459667,-0.0298742855637915,-0.0157296555964452,0.0100996020885236,0.00271188526589716,-0.00774642455607477,-0.017418389804244,0.0174113214902445,0.00266307934858157
"2174",-0.0301025244679525,-0.0216113554222853,-0.0340357023653962,-0.0307783139121482,0.0030154822479358,0.0040106976832841,-0.019584754014182,-0.0206409083002371,0.006247690940824,-0.0166002437314864
"2175",-0.0421068263941223,-0.0268907325722504,-0.0352347660945919,-0.0436641014417188,-0.000316451744231117,0.00167207005620318,-0.0466999760739935,-0.0453757449285994,-0.00539906430484294,-0.0249831944517125
"2176",-0.0117679032975058,0.00616814436375002,0.00608691690119811,0.0127713244233978,-0.0160650187430929,-0.00547174574871612,-0.02520185984803,0.00701321261114485,-0.0123947798099592,0.00415521063827451
"2177",0.0383939858634177,0.0166746739711499,0.0397579860390878,0.0331022258117681,-0.0193035934920132,-0.00615394048538109,0.0249818406112561,0.0201183932194857,-0.0136497429956122,-0.00620695348291322
"2178",0.0247350465552016,0.0108540808666475,0.0182877027936712,0.0442479018906528,0.000574212897365811,-0.000563213498712356,0.0201218379694028,0.0199746815593678,0.000557304737759834,0.0360860590358638
"2179",0.0000501038309095314,-0.00238619178392141,0.00489790174274685,-0.0128582409218236,0.00295083773469096,0.000187492538685996,-0.00111105194387973,-0.0101634722057422,0.00900393551460321,0.0261219592799926
"2180",-0.00807885603954539,-0.00454430161478014,-0.0154346983150987,0.00177613358915085,-0.00768251099650241,-0.00168925364598793,-0.0198860799996985,-0.0120210201872664,0.00110398347113105,0.0241513737615482
"2181",-0.0298479459000403,-0.0285920466648837,-0.0453794687968112,-0.0387113061237917,0.0072055354053,0.00449184288645488,-0.0190124181898196,-0.0263625830073452,0.00349197757765118,-0.0331421357263799
"2182",0.0189811988052271,0.0140984356217277,0.018150365516362,0.0144481359869144,-0.00860439458588413,-0.00271878740409792,0.0107029979651372,0.0179639526698487,-0.00531130051221518,0.00856963182897941
"2183",0.00071641063132355,0.00146346992628299,0.00764009450204073,0.00393942884118426,0.00487677006175069,0.00244454219690526,0.00200313560008469,-0.00306884462326562,-0.00718106222110859,0.00653585802039114
"2184",-0.0151368231199519,-0.0211884106169564,-0.0320135568448837,-0.0298823226721946,0.00913028065937471,0.00309425734996704,-0.0189943106956684,-0.0218061013364784,-0.00324553053581345,-0.012337627793219
"2185",0.0251310912902569,0.0291118165422231,0.0234987775622384,0.0317360936634954,-0.0147537099420516,-0.00439372429936735,0.0151404974361522,0.0251773081771289,0.000279086431837161,0.00723212063576195
"2186",-0.0133716454282371,-0.00531935784111026,-0.00170065274581277,-0.00512655933449724,0.00479862803473896,0.000374879037473574,-0.0121899418268672,-0.0138147147952223,-0.0129278277416619,-0.0130548529148178
"2187",0.00544156262911533,0.0094798205853186,-0.000851740204090179,0.0103062573586932,-0.00675173399685058,-0.00225228654274301,0.00116149784961506,0.00985747288358785,0.00235560168724014,0.00859783403115144
"2188",0.00454438046168337,-0.000963066709138483,0.000852466283896902,0.00390039056166325,0.00629988828422956,0.00263445330839929,0.0163860885456644,0.0020548989709066,-0.00206799216209796,-0.00131145753062911
"2189",-0.0037105049876075,-0.0106049684014617,-0.00255538274261879,-0.00149452199923295,0.00156567740038782,0.000938183932521541,-0.000570671469845574,-0.002819571775177,0.000565156346452156,-0.0124754099800847
"2190",0.012499369297075,0.00682090908052579,0.00768576513797536,0.00957790702796268,-0.0191645710089287,-0.00787411399167326,0.00842294010795031,0.00385592362773757,-0.00301260588389562,0.00332449124458023
"2191",0.00866662728651213,0.0164531070514404,0.00847446183378975,0.0243107785021048,-0.00377325234764414,-0.000283561079739258,0.0128819314148116,0.00717038770591616,0.0133144095691329,0.0165673099142225
"2192",-0.00224797966195467,0.00285643353674914,-0.000840288322131122,-0.00231535628286483,0.0122052282158893,0.00831673274208833,0.0097836515206422,0.0010169657932102,0.0102507317165359,-0.00651901687994838
"2193",-0.0163414115292977,-0.0256350318043432,-0.0319596166888683,-0.0185670029204447,0.0153846987255479,0.00468687746570273,-0.00332181274646248,-0.00787739730665116,0.00737934665144002,-0.0150917261893305
"2194",0.00516758087237168,-0.00219275421250176,0.00608172332700629,-0.00177350832582523,-0.0162982516125469,-0.00569087708910354,0.00874837733173917,0.00438235816157717,-0.0062265360885132,0.0113257646300211
"2195",-0.0129796597768439,-0.0302730849831385,-0.01468042150229,-0.0186556164241161,0.0139043103026602,0.0049725221919259,-0.0132157015223162,-0.0148869017707549,-0.00681837286297216,-0.0059289081563676
"2196",-0.00159869560466663,-0.00377657706039769,0,-0.015992661229502,-0.0000825368841204099,-0.00112002673045297,0.00460404017469385,-0.00338751437014706,0.00398923829678788,-0.00795224601006539
"2197",-0.00361588184986206,-0.00404333986147487,-0.00701156528400093,-0.00429326506220007,0.00681610075512418,0.00149538904006086,-0.00916561148607631,0.00967328667112466,0.0209757621421571,0.00601201054571754
"2198",-0.000259014797913237,0.00659719977007822,0.0247131606494519,-0.00215587113727589,-0.00864574330677281,-0.00261324625703452,0.00503666221407406,0.0137237309931681,-0.00615440322480598,0.00597601393501157
"2199",-0.0250973008783402,-0.0186537796903842,-0.0241171496556061,-0.021296337363566,0.0171137565384536,0.00570784623307263,-0.0180181949179805,-0.0153260351146324,-0.0126582280786489,-0.0138613336739144
"2200",0.000585048916816655,0.00436670164217223,-0.012356496326029,0.00473044105829312,0.00283115012328228,0.0034420063099514,0.00702426338515649,0.00337254261630027,-0.00405824578598513,0.00669341801839107
"2201",0.0186583474998208,0.0179027068231292,0.021447884112662,0.0288762018725295,-0.00346867525600847,0.000185907994777912,0.00996402659734974,0.0170630626239185,-0.010372309398806,0.00731379861976911
"2202",0.00260916153351332,0.000251505808943175,0.006998939267018,0.00549132569941646,0.00426663801999716,0.000779697183793004,0.00465116695445933,0.00152488393867567,-0.00121652628470403,-0.00660057038275963
"2203",0.0149378207705093,0.0198440364975281,0.012163352156787,0.0266987644453303,0.00605755573433431,0.00482454957069289,0.00869853588891689,0.0114213764143247,0.0211748799444895,0.00664442739342297
"2204",0.0177948322122352,0.0189656035048729,0.0248926627114168,0.0215722796735773,-0.013567583725804,-0.00553957838645569,0.0179412678528841,0.0225847699224131,-0.00201854302263582,0.0132014125057576
"2205",-0.00342613721428631,0.00459282704537478,-0.00837509692408145,-0.00173554487239747,0.00431336058520682,0.00204229171830339,-0.0024593914604627,-0.00318991157711679,0.0100211825876946,0.0195439748149826
"2206",0.00819055532945612,0.00962434803408674,0.0160472086149521,0.0266589463382387,-0.00332275047684638,-0.00250158937547895,0.00972492588394513,0,-0.0014564354500598,-0.00191690668555067
"2207",0.00902663676277582,0.0088181829532068,0.00332496700732765,0.0107253136512759,-0.00837412442901864,-0.00260064083200962,0.00827449898120824,0.00960104644414228,-0.00510481326631207,0.00448137263945814
"2208",0.000596448659801574,0.000944946705688343,0.00248551749966164,0.00363042790800749,0.0026235320926995,0.000558547241255036,-0.00107612284993697,-0.00414525760806339,0.015851237088613,0.00446151072916767
"2209",0.0009435127187849,-0.00354018454965177,0.00165286589228497,-0.0075128327112407,0.00760546599800827,0.00335059655544168,0.00538713699045101,-0.0019589691216797,0.00396856668254975,-0.0158629878376184
"2210",-0.00630206498017638,-0.0106584760109691,-0.0107259559141054,-0.0162599511169413,0.00170460570492215,0.000927712667972314,-0.00736759688064237,-0.00981335339349521,0.00494118237249452,-0.00644743147882887
"2211",-0.00479421143515124,0.00526692556924924,-0.0116764116373593,0.00769453363641426,0.00875047415132313,0.00546806778535758,-0.00647792515039847,0.00941515005518934,0.01743247794178,0.00259568152702783
"2212",0.015354742052156,0.0126218631702451,0.0253164583103582,0.0243211776126802,-0.00489942691628897,-0.00341040828980543,0.0114100520151856,0.0130092884276907,-0.00456899226024055,-0.00258896140772769
"2213",0.00454670059225593,-0.0018815566175322,0.00493828105422822,0.000828333583343888,0.000322746658708128,-0.000832573565499262,0.00805787545791081,0.00314991169054535,-0.00706154994208186,0.000648920381757012
"2214",0.000491688578591942,-0.00376977491582742,-0.0049140142706553,-0.0102067450571826,-0.0027435667291541,-0.000462483055415852,0.0118571541951811,0.000966251688571784,-0.004178158132779,-0.0181582545830651
"2215",-0.00127815154671684,-0.00307475609896635,-0.00576136892641199,-0.000279111380814046,-0.00614922590773226,-0.00342681984125925,0.00118509563193325,-0.00120660857640242,0.0063382076326961,0.00198147886929001
"2216",-0.00620358254732978,-0.0045079436896498,0.0132451116725201,-0.0144966455571452,0.00993242557268892,0.00343860331532642,-0.00355115732858147,-0.00507391033099835,-0.00887075289086969,-0.00856956398348829
"2217",0.0168936261582782,0.0102479518207177,0.0122546918407038,0.0206507384256751,0.00169278216578683,0.00101836407535782,0.0109543999874355,0.0179703353385006,-0.000358014847632204,0.00332449124458023
"2218",0.010961613067028,0.00825666974938177,0.00968542589443899,0.00582040055407629,-0.00853055536889991,-0.00564320290718379,-0.00913838914602538,0.0023851721381114,-0.0017011549520789,-0.00596420155884292
"2219",-0.00245760192738509,-0.00491342788961879,-0.000799314937497297,-0.00909350870592451,0.0066560062715697,0.00260484302387187,-0.000131602649806384,-0.00380756799983495,-0.000627802690582935,-0.00266663025528879
"2220",-0.00193243948442579,-0.00940492399088488,-0.00800004385457054,-0.0114015922304593,0.00249935736048457,0.00250560757541729,-0.00250352713098967,-0.000955601716360333,0.00224356097998735,-0.00467914912177814
"2221",0.0113746063533593,0.0073578639545071,0.00967743774664309,-0.011533087794652,-0.00402143861826521,-0.0051837830904834,0.00383072258254957,0,-0.00805874820916908,0.0167897693851011
"2222",-0.000574354892483586,-0.00424109131909944,-0.0111823613380636,-0.00939082062869145,-0.015909074753798,-0.00614111121100147,-0.00105267814330279,-0.00645638602564924,-0.00956849620480682,-0.00594450458779516
"2223",-0.00430960894183186,-0.000709945029986114,-0.00484638326815445,0.00172357886617869,0.00754986549011316,0.00196613887788333,-0.00724560564716403,-0.00216601793866711,-0.00382790736576821,0.00996670947658385
"2224",0.0118310091985399,0.0113664304890186,0.00730522040550463,0.0197877888973343,-0.00459558762175294,-0.00287298363082233,0.0221602520209159,0.00554743413131531,-0.00649594675674436,-0.00526308626300498
"2225",0.00289924461234503,-0.00210726047334853,-0.000805733973956113,0.0132170073990361,-0.00820001753335531,-0.00262804707308861,-0.00986620328428389,-0.0040775181990258,-0.0148263473552389,0.0178571708144006
"2226",-0.0030333549887388,-0.00680426867230788,-0.00483880658808011,-0.00804885117527776,0.00115731571555489,-0.00103482349351924,-0.00432642304723907,-0.0144507643142596,-0.00944103544285746,-0.0168941229624917
"2227",-0.000998085146887928,-0.00307101586063241,0.0072932923908382,0.00167872941671043,-0.00264222459042252,-0.000659618742285262,0.00289684117954248,0.00171032848640085,-0.00311410773696219,-0.0079312219733344
"2228",-0.000523490826623285,-0.00545035092978752,-0.00241335659135822,-0.0139663617888904,-0.0146559275329994,-0.00678662622616921,-0.0286238152847116,-0.0124419409016485,-0.0145778210391692,-0.0059960575746596
"2229",-0.00933152743762355,-0.0104837911636864,-0.00403224745385977,-0.0249291863555748,-0.00563050035804202,-0.0017082991657914,-0.0135173277050903,-0.0249505713333704,0.00288188286036273,-0.00871308670317672
"2230",0.00230669647786619,-0.00433413142644845,0.010526199908055,-0.00435783553017388,0.00295781004204976,0.00190117901410214,0.00918062839820233,0,-0.00210729881020499,-0.00202843934733932
"2231",-0.00393146312044157,0.00507867774012283,0.00400648728301323,0.00204257074393954,-0.00210639376559407,-0.000474052613679499,0.0012219256973629,0.00810765832959381,-0.00335955077750061,-0.0101626021929274
"2232",-0.0139599243477254,-0.0153995967804665,-0.00957705532723974,-0.00961001461360822,0.00481312845176318,0.000569276369193572,-0.00718745772537777,-0.00804245286959537,0.000192584027880471,-0.0143737315317003
"2233",-0.0112283402304991,-0.00855339224430729,-0.00483473250905087,-0.0138193731768523,0.00571388219348834,0.00379510447613352,-0.0105175111681257,-0.00481372632248445,-0.00279248922084718,-0.00763885608064085
"2234",0.0152070123646719,0.0125710588200392,0.00971663957050062,0.0193798527032654,-0.000918991027511695,0.00132341624561017,0.0117337525803833,0.0132381389797933,0.00144844537366651,0.00489846340708389
"2235",-0.000729468650744525,0.00316465763308482,0.00240576740476062,-0.00292463702156642,0.00167269206712328,-0.000283144993562634,0.000545909213626627,0.0047735132771074,-0.0132099413095164,-0.0153202689780357
"2236",0.015866072395877,0.0101916668945365,0.00480003066339418,0.0108534283746637,0.00208765416197454,-0.000472128127406823,0.0106366269366396,0.0072522196254845,0.000879460655831998,0.00424322340568328
"2237",-0.000862318711467136,0.00576512495106041,0,0.00899616762993283,0.00666531569364559,0.00217251529494078,0.00283377040361832,0.00571004491167848,0.0110319047154153,0
"2238",0.00364412349233234,-0.00740388264135261,0.00477684064272488,0.0100660863692164,-0.00306245716316689,-0.00131979864432596,0.0102258323772118,0.00444341467728049,-0.00453845122708474,-0.00140843151233594
"2239",-0.00114689211160235,-0.00697792332782676,-0.00475413091693999,-0.00939648461624187,0.0030718646169674,0.00132154281474128,0.00173180222594493,-0.0105676759174597,-0.00805115949369128,0.0077574441065984
"2240",0.00133944522387752,-0.00169622043610351,0.00477684064272488,0.00517393446730519,-0.0000826265177638064,0.000942726586306675,-0.00491957794184184,-0.000745382379443327,0.00664971627909816,0.0160951672652541
"2241",-0.000143135196755573,0.00582529550307109,-0.0063389776832331,-0.00772084223817004,0.00231723893681757,0.000564874319536557,0.00334025128417736,0.000248745283969898,-0.00466293948585716,-0.00137739162486072
"2242",0.00114652099238932,0.00482620609577777,-0.0047848064408732,-0.0219020872847689,-0.000990954494104024,0.00103525527290382,0.00799039992712269,-0.00472164771042072,-0.0118094769842814,-0.0151724188841127
"2243",-0.00415153031148319,0,-0.00801295277790293,0.0014732213617985,0.00396814805563506,0.000376351628373461,-0.00634141964613666,0.000499195182228629,0.00661726419753084,-0.00630257884926444
"2244",0.00953556357801699,0.00696454556821946,0.0153474294521774,0.00764940943158554,0.0135071894945775,0.0053182166870227,0.0123652223713062,0.0187173813067565,0.00353219198454058,0.0112756100009341
"2245",-0.0102049821160304,-0.0114477535283278,-0.00795525663518337,-0.0119710986665251,0.000325729480815218,-0.00280875751033205,-0.0189127336791739,-0.0142086974032248,-0.015545532025279,-0.0209059238447552
"2246",-0.0140027887819353,-0.00506623194042055,-0.00962313503581946,-0.00561442902022036,-0.0271831544686735,-0.0105166202769876,-0.0147255602660076,-0.00670969425222101,0.0106266757249642,0.0113878176129558
"2247",0.0195029512921314,0.00994175184978219,0.00566789113153932,0.00683500231543133,0.00878451997687213,0.00370066186591878,0.0167121395502454,0.0085062639723239,0.0222090699251363,-0.0014074403706511
"2248",-0.00605854417289475,-0.00672273130903589,-0.00241554042922454,-0.0165289640238293,0.00970304785944931,0.00321485267288635,-0.00267284360342435,-0.00868267037304604,-0.0129782641697249,-0.0288936282311872
"2249",-0.00671956285939346,-0.0157117590648399,-0.0129134768956609,-0.0111042783174142,0.000492409482168332,0.000565525882975093,-0.00241163201042938,-0.0102601105820607,0.00165577094878278,-0.00507975678233286
"2250",-0.007779706264891,-0.00221032736993865,-0.0114472755230348,-0.00819430312706737,-0.00106709786211223,0.00150694550984709,-0.00617859346893457,-0.002781426450985,-0.00194473947665263,0.000729459707354385
"2251",0.00258113266424886,-0.00319962341704272,0.00909844990246667,-0.0067320504848265,0.00131517680684823,-0.00216332102712902,-0.00567661773944217,-0.00329616780794695,-0.000876812167544982,-0.00364433985582713
"2252",-0.0193811795916975,-0.0170368873143667,-0.0155737744561757,-0.0280346178077143,0.0157582088224144,0.00801157176546607,-0.00462129747296547,-0.0167896046901449,0.00546073119081236,-0.0102415653600367
"2253",0.00505244218358869,-0.00150698527730619,0.00915894236859827,0.0161649319302555,-0.0129280730628901,-0.00738688401675136,0.00314057564160963,0.0049160265520547,-0.0128018619648738,-0.00665179463204035
"2254",0.0104978006107674,0.00905619271459046,-0.00412540217511081,0.0152838834775628,-0.00589396874160775,-0.00254317934870518,0.0110261676370704,0.00334698391447064,-0.00265255916443108,-0.00223211243083221
"2255",0.0146319978596436,0.0184493524078102,0.024855107411915,0.0196622023293955,-0.00214104719855535,-0.00264417741089795,0.0196582848765208,0.0207850725964656,0.0121158691523602,-0.00447421180545382
"2256",-0.0152381411597808,-0.0141981017787258,-0.00970084189030818,-0.0129559140167667,0.0113055624063736,0.00416627914709977,-0.00488590928505539,-0.0145802350129201,-0.0218978102189781,-0.0104869787599111
"2257",-0.0178149174270763,-0.0124163341696536,-0.0122450207233091,-0.00335758431435418,0.0055487386526023,0.00358338452795248,-0.0127386801985058,-0.00282349276230665,0.015323393034826,0.00454210752137274
"2258",0.00824902522675597,0.00475451402405369,0.00316361646454966,0.00780737321379976,-0.000243696882155864,0.000469791192718505,0.00510731388184515,0.00360395559204485,0.0108780967181683,-0.00452157006397669
"2259",0.00907440128061388,0.00729919866685269,0.0074689317399379,0.00802470176840697,-0.00722361764016954,-0.00281759808656501,0.00414560864217872,0.00487304655228082,-0.00523510411565486,-0.0045420296094798
"2260",0.0123833117434491,0.0194901785268011,0.0107083624330304,0.0140843723898472,-0.00752219229070306,-0.00226039602410966,0.0113200258205204,0.00995406085308681,-0.00292372085641046,0.0182510150888562
"2261",-0.00165056072080383,0.00147062126520092,-0.0122252072842475,-0.00362303012550436,0.00572949698501479,0.00183409558956349,0.000266491019621951,0.00151622355868097,0.0072329685706769,0
"2262",-0.00228474201345008,-0.0041604137166259,0.000825249328729072,-0.00696963015543439,0.00295479025769052,0.000188520409978965,0.00293338114284558,-0.00656054408575324,-0.00756919919740318,-0.0141898071176862
"2263",0.0106716523677479,0.00884724374264922,0.0148392573641778,0.000915313842738019,-0.0166135065450228,-0.00528344642666234,0.0102366167817154,0.0104137844802918,-0.000684462716861178,0.0166667524346811
"2264",-0.00708769684279842,-0.00803881010150609,-0.005686529915084,-0.0155487537949011,-0.000998603487003535,0.000379448257469939,-0.00447422966599476,-0.00703846893517734,-0.00763208437276164,-0.00968705542198245
"2265",-0.0100034928094693,-0.0149805518373126,-0.00980400632431733,-0.00309704813950518,0.00449845854002828,0.0011379026445042,-0.00753461964716984,-0.00962059123286918,0.000394409394486317,0.00526712378627625
"2266",-0.0139794726430926,-0.0149588013203923,-0.0156763964259642,-0.0273376272515576,0.00721492573762816,0.00426156901162811,-0.00972303753031234,-0.00894701082068339,0.0140942244637712,-0.00748492787745059
"2267",0.0016914466130602,-0.00632754317735729,0.012573350275406,0.00223584963831303,-0.00403458374731414,-0.000282794702954892,0.0164090245417621,0.00154805615773457,0.00281855382270924,-0.0098039421145949
"2268",-0.0126143144658164,-0.016811090350012,-0.0173841540556964,-0.0191204610347214,0.013475694125715,0.0060369459643328,-0.00330863002524873,-0.0100439872193487,0.0144407637138981,-0.0159939228439159
"2269",-0.0239912763087226,-0.0181346116016324,-0.0151642964029811,-0.0308643141694728,0.00179458935745025,0.00215700221457005,-0.0223046770776557,-0.0228927783025503,0.0141397155658682,-0.00464405853976857
"2270",-0.0109767425940933,-0.0100264696199635,-0.0213859417747193,-0.0107275268981515,0.00447855907081385,0.00252627181864118,-0.0118139178233874,-0.0135782234734825,-0.0044277154135145,-0.00466564641415823
"2271",0.000990112894379225,0.00346499291800328,0.00699326489895169,-0.000338884428674024,-0.0109437172812746,-0.00317342341142446,0.00398487823984062,0.00377858186543945,-0.00889479560938689,-0.027343700059397
"2272",0.00806827980883429,0.00796818429712687,-0.00520835420257781,0.00203395859251621,0.0144250089897719,0.00449395576510181,-0.00698064253259423,0.00430224010495972,-0.00506013948940498,-0.00642569783124736
"2273",-0.0249407310819555,-0.0171277857286932,-0.00872614070850952,-0.0104871636637704,0.00985698668260304,0.00391509476862684,-0.0151619124003004,-0.0109771020153471,0.00489398334990865,-0.00565877484512667
"2274",0.0164167628328937,0.0128685218667792,0.0123240821351696,0.0129915493698911,-0.00936078370168902,-0.00204300034016403,-0.00139947806276286,0.00893345500086062,-0.0162338042758421,0.00243899091980437
"2275",-0.0214660146857475,-0.0367920874174253,-0.0278260738933502,-0.0394869655499992,0.0155873984815877,0.00465161444556927,-0.0113524596987723,-0.0300511378591172,0.0102893130544353,-0.0210869089061161
"2276",0.00133103911435173,0.00906861380937118,0.00805007348572229,0.0147574484241064,-0.00310153559319692,-0.00129665648520438,0.00297730830254439,0.00553250482299705,-0.000960789758632008,-0.00828489181420122
"2277",-0.0128150121177718,-0.0206972778827144,-0.0381545779625333,-0.0218143451402258,0.0105298621980734,0.00491459266985284,-0.02657300500307,-0.0220080403632341,0.0133679549903456,-0.0075187801837816
"2278",0.00560207935926615,0.010845611173909,-0.00368993628137604,0.00389383587940229,-0.0067889623336318,-0.00249121736282631,0.00667955176090795,0.00450063644800669,0.0011387965890064,0.0134680023834841
"2279",0.0205152520995848,0.0264097376108798,0.0453704908289116,0.0342030708792158,-0.00381496526071623,-0.00221992785254677,0.0276936574470019,0.0229626059690105,-0.00464497117537155,0.0299002652026497
"2280",-0.0151166144776743,-0.0134012679001075,-0.0212578115305446,-0.0170473449853906,0.00542520522818091,0.0033373711746616,-0.00982459091149368,-0.00848612171427643,0.0102857333333333,-0.021774146157322
"2281",0.0136429690277569,0.0214613950680889,0.0135747647598483,0.014568015310507,0.000476013157693522,0.000739101676612508,0.0214032617680757,0.0168415983012167,0.0114064760292898,0.0197856396611851
"2282",-0.0108829801731624,-0.0085105676099414,0.000892844618620936,-0.00341866656142131,-0.000237822552699107,0.000738626350892835,-0.0155424961550202,-0.00705945242821859,0.00372822253958227,0.0121261125018888
"2283",0.00520906531207355,0.00214619521791448,0.0017840722363236,0.0157803703031651,0.001428106685186,0.00129179060579898,-0.00662558482051412,0.00710964261201985,-0.0106788093475939,0.0111821204449172
"2284",0.0243774057562294,0.0160597953897141,0.0240427434027635,0.0324215457415347,0.00847657194529949,0.0053435539431923,0.0217115792867546,0.0285094333786804,0.00384828229915257,0.00947862482423667
"2285",-0.000361439333254499,-0.00158064654247581,-0.00608689498195458,-0.00948648241082595,-0.00306163341080412,-0.00230336997667802,0.000138867234821483,0.00712769027501547,0.0102852363801376,-0.0187792482003014
"2286",-0.0180221781860751,-0.0274404764357168,-0.0104986820853086,-0.0323645846230598,0.0185523033616741,0.00708365217264717,-0.0105540876287016,-0.0212320839764264,0.000370134186854276,-0.0175439474833902
"2287",0.0059949453427961,0.015192567138214,-0.0123784433913752,0.0283276869929294,-0.00829343105372315,-0.00109623966110606,0.00491227884876477,0.0182111300801779,0.010731834979437,0.0251624127265246
"2288",0.00156822668982115,0.00133620858755457,-0.00268596946170296,0.00763366076580785,0.0048456346389778,0.00237785070407437,0.00111739214637341,0.00236705559139549,0.0120823798627001,-0.00158359108553852
"2289",-0.0190499034220524,-0.0152121284553914,-0.0170555893449515,-0.0115285148498931,0.00116679416411869,0.00127766888856873,-0.0224611651209837,-0.0170557826092083,0.0158270778692231,-0.00634416643820135
"2290",-0.0134611747952191,-0.0235773740163043,-0.00182633540900634,-0.0136619979610042,0.0215195283931577,0.00747130124847284,-0.02939890005757,-0.0149489710512868,0.01344375,-0.00478852442938482
"2291",0.000053789184865316,-0.00888160206942978,-0.0192132262889751,-0.0138513449140438,0.00106458540390975,0.000180640837911694,-0.0161740392752862,-0.00406555033788447,-0.00219625753850028,-0.0256615684840983
"2292",-0.00086268030872505,0.0042005187635088,-0.0177238847076868,0.00411092975487137,0.00881283909378627,0.00298361298303207,0.0052309043105585,0.000272215020091338,0.00774781638056332,0.0016460680853132
"2293",-0.0130082588491816,-0.0142218649970429,-0.0199430745729247,-0.0167177811704071,0.00700311544827925,0.00459843195403153,-0.014719219522644,-0.00843295387347698,0.0401887038283129,0.0123253916243458
"2294",0.0206170475301601,0.0195190961530083,0.00872099197477882,0.0173490150216573,-0.0166016930305537,-0.00762827423664814,0.0129772275469451,0.0150889202895204,-0.00587936344497497,0.0146104412805887
"2295",0.0168782080391958,0.016092978321318,0.0365032927791613,0.022169216095457,-0.0105702527643995,-0.00298440525912136,0.0192164825091941,0.0202705364565243,-0.0303312265095367,-0.0112000939303752
"2296",0.0163348445346283,0.0207539587770582,0.00834111563434825,0.0196861201209459,-0.0061487933695511,-0.00244910150463129,0.00906170066592171,0.0127150789808066,0.00618633805488367,0.0210357295389787
"2297",-0.00409594528016533,-0.00588546918854627,0,-0.00588986755344045,0.0122962064625638,0.0046375064453168,0.00955957332960944,-0.00392328412923793,0.0243331999220679,-0.00554667519181595
"2298",-0.000468349310332239,-0.00188379311898523,-0.00459574733715773,-0.00460837064530872,0.000840301208675731,0,0.00215220339200584,0.00787792497527962,-0.00600218948345443,-0.00876506550734024
"2299",0.0144790438530806,0.00727973763898415,0.0166207177620281,0.0248017214042575,-0.000534442699552828,-0.000995437769243268,0.0115963159587382,0.0104220962406121,-0.0177751655421812,0.015273351601643
"2300",-0.0126296861398921,-0.0173986379347831,-0.0163489858819882,-0.0212972170268891,0.00404780327379828,0.00199278031352645,-0.00240589725400531,-0.0167615175265198,0.0149796781536007,-0.0134600760332335
"2301",0.00457575287509493,-0.00435832509392475,0.0101570803739723,-0.00230802002794883,-0.00197745215687462,0,0.000425374833350256,0.00550778703565435,0.00332707726218162,0.0128411642829631
"2302",0.0121118315310353,0.0139535360909917,0.011882956175705,0.00330485091510857,0.00358139698370952,0.00298402376434348,0.0181512067666194,0.00834604471119005,0.00263580475609393,-0.000792463724620274
"2303",-0.00230146187493807,-0.00296809799041364,-0.000903232294344969,-0.00988156863705114,-0.00964429589239379,-0.00486801855999131,-0.00306444561157815,-0.00646618219153616,-0.00686903844757536,-0.00158593958574915
"2304",-0.00784253395563794,-0.00460103278393553,-0.015370758757926,0.00864941628345184,0.00437106717939373,0.00163080815955396,-0.00167635024383539,-0.00104159502418,0.0130646228924549,0.012708406021543
"2305",0.023507105225935,0.0274607560492541,0.024793390068609,0.0356200521485561,-0.0176088444580764,-0.00781613171770812,0.026028681948278,0.0242377715128743,-0.00733312548325293,0.00078430302575816
"2306",0.00449236427116295,0.00238174123054735,0.0143370080727001,0.0133757706650199,0.00412707726842987,-0.00173466357256769,0.00763764276775269,0.00585221118897605,0.00772695103320764,0.00548589929572096
"2307",0.00391969606268416,0.00844753604705795,0.00706703871714698,0.0113136277974701,0.00364461901384883,0.001188805487641,0.00500810976232424,0.00455357534176559,0.0172733653522075,0.00545596840250417
"2308",0.00325352827559788,0.00523569941638291,0.0105263823393358,0.0198881246013987,-0.00641296096851873,-0.00337955084912478,0.00269377268827431,0.00302232226114718,-0.00157377615570831,0.0193798199127144
"2309",0.000798200082179346,0,-0.01041673183729,-0.00152329973931409,-0.000311008984338224,-0.00201598133431447,0.00188030644533854,-0.0057750335812744,0.00497758416311944,0.0182510150888562
"2310",-0.0109179436968657,-0.0106770492534617,-0.00964905949741102,-0.0170889450070237,0.0110454294864115,0.00578496550784702,-0.010322998189103,-0.00303008378833425,-0.00462272580999457,-0.0134429144816003
"2311",0.00493992725281278,0.00552763847740656,-0.000885894570130108,0.00620930999527802,-0.00607817913801534,-0.00392581145614002,0.00406394684638345,0.000253458527296191,-0.00829324915751783,0.0151400727276354
"2312",0.000802321015206608,-0.000523552039363051,-0.00443249100959708,0.0015426378486425,-0.00410221400066557,-0.00357459696451656,-0.00256355377287276,0.00177252192453037,0.0160561796946617,-0.00149140393515124
"2313",0.0161371880754044,0.026715469154253,0.026714170019621,0.0209489150629711,-0.0101041927201015,-0.00285162540545703,0.0236710499324246,0.0245199563898735,-0.0172016131687243,0.00373407885778065
"2314",-0.00128233071757877,-0.00280606434153063,0.00433640600876317,-0.00603512584903632,0.0031408939912414,0.000738110196932817,-0.00132131920098766,-0.00197399611206794,-0.0128967502588812,-0.00892852630190855
"2315",-0.00162975064997573,-0.00946529093968762,-0.0129532115246835,-0.0142682166526533,0.000939091729644348,-0.000184230924429429,-0.000264735592469978,-0.00296703040725099,0.000763519111813382,-0.00825829985097226
"2316",0.00578714215417242,0.0103304464742424,0.00174973311427484,0.0200183521651829,0.00297163775154052,0.00525529675710579,0.0127052864659718,0.0126459872634757,0.0222956682120692,0.0174110485764289
"2317",0.00634401029911413,0.00741322068252459,0.00349335379174032,0.022041123460008,0.00413188795874553,0.00110070779579985,0.0139832578518222,0.0173847378339598,-0.00381457015721265,0.0111607918898995
"2318",0.00392994039437733,-0.000253753198956264,-0.00348119275383385,0.00531757228984886,0.00209642127858412,0.00174041248049983,-0.00386660708796527,-0.00166686354281786,-0.00274697417997938,-0.000735900819623936
"2319",0.00141886594527318,-0.00482241880020684,0.00436679832891995,0.00205701008839254,-0.00767041790618361,-0.00283497602310012,-0.00646908405285396,-0.00121014972341293,-0.00701171935696865,0.00294554370651778
"2320",-0.000537524134409884,-0.00535564977128289,0.00608705929215869,-0.00234589544870178,-0.000234438949827331,-0.00210941044274515,0.000260749004829197,-0.000727033370522268,0.00294215705230449,0.00734219461659547
"2321",-0.00659944774801591,-0.00820505812488481,-0.0129646611046494,-0.0170488329956437,0.0113247823483917,0.00459521704061339,-0.00704837022671378,-0.0106692756297103,-0.0226300984432167,-0.0211371111512028
"2322",-0.000442988360693453,-0.00723891657201914,-0.00612962975613307,-0.00239236015000344,0.000385874606853687,-0.00100629081369386,0.000796111655082532,-0.00661732237186363,-0.00240115768457971,-0.0059567318472874
"2323",0.000590884266200797,0.00416663092492775,0.0149780264359161,0.00329725602833175,0.00131263438737994,0.00146517102237298,0.00768920564924058,0.00320684056697806,0.00232094898442448,0.00299621356440394
"2324",0.00924997358830737,0.0121887091853172,0.0104166615408874,0.0137435865901403,0.0104846187247098,0.00676744866616974,0.0198654792019219,0.0150029334069515,0.0185249059781287,-0.00224052417919829
"2325",0.00438783704910795,0.0107609314747694,-0.00343651720555638,0.0103155906073533,-0.0105287622509055,-0.00136238020314439,-0.00154761133506132,0.00823841437891026,-0.0139778037390064,-0.00374246393872524
"2326",-0.0024269307049829,-0.00861857258968812,-0.0163793155004549,-0.000875219694928764,0.0070941072454358,0.00363806256883548,0.00594279329504288,-0.00360502063765245,0.00461145182940137,-0.00150268636214512
"2327",0.00681180747556165,-0.00869338156286892,-0.0245398440632472,-0.00291975128265765,0.00260843259016852,-0.000290483184007484,0.00064254778901307,-0.0089242357093765,-0.00603535367252084,-0.0173061642997535
"2328",-0.00323803402277223,0.00128971040988857,0,-0.0120058835812503,0.00061207420763254,0.00118039506437673,-0.0014121871240016,-0.00292023249986961,-0.00667064055417776,-0.0137825107354482
"2329",-0.00998773641174455,-0.0190623941367132,-0.0215633331659053,-0.019561310311197,0.0109362204568799,0.0039903721376422,-0.00565526396194105,-0.00610231064999578,0.0130004474730874,-0.00232932034986943
"2330",0.0109211419795587,0.0152311551446249,0.0165288688744074,0.0120918452589724,-0.00726227349877717,-0.00216814426703915,0.00245595056326886,0.00982320430558037,-0.00611934366413924,0.0108950335716682
"2331",-0.0119657971565379,-0.016813202558575,-0.0054199058439891,-0.0200119204188894,0.0123448456708573,0.00516015514560464,-0.0054158094519976,-0.00851177171497419,0.0142808189792916,-0.00307932878634831
"2332",0.0026965364056275,0.0176270394599833,0.0290642753691073,0.017372779294851,-0.00632322940606433,-0.00153107819709242,0.00570438792493944,0.012999832746007,-0.00151758703720095,0.0239382940858939
"2333",-0.00234694764647436,0.00180964810914697,-0.00617813088144603,0.0128819225825134,-0.00128758738340284,-0.000180524135330984,-0.00128899550574557,0.00411618400205316,0.0135100819049228,0.00754137452184356
"2334",0.00931277182504409,0.011354719688851,0.0230905990477415,0.0153801834176939,-0.0069025743467418,-0.00396933649107301,0.00684150482133883,0.00795775207867666,0.000166658336804515,0.02170659899314
"2335",0.0101008433278589,0.0137791600663111,0.0277777641090329,0.0177687312028088,0.00351346982997303,0.000724927944697695,-0.00230782014719533,0.00885151955048458,-0.0106622737860324,0.00512828594201653
"2336",0.0000481865228223466,0.00125851814157829,0.00422302794820095,-0.00486536980740704,-0.00479489924357179,-0.00235337968813643,-0.00642497782044815,-0.00545398582834633,-0.0139765600903401,-0.0080175326796712
"2337",-0.00110572932390285,-0.00175960762294358,-0.00925165986436838,-0.00575226418505748,0.00856550204803219,0.00299403975080104,0.0065958565101889,-0.00238433215927791,0.00691654848504375,-0.00367379462428574
"2338",0.00702665397598246,0.00906558353217979,0.00764012257303648,0.00462828903607626,-0.00432238097429805,-0.000995332224577816,0.00424001534595919,0.00693119625407879,-0.0015264586419006,0.00442479420991582
"2339",0.00315423044852325,0.0197154314983372,0.015164410109052,0.0152605196927096,-0.00312239665316161,-0.00162971493694009,0.00102348690992793,0.00593397885701119,0.0156276883918411,0.0212922283683834
"2340",0.000952922328843142,-0.00244731531317732,0.00580886795522684,-0.0045376563552304,-0.0110004736112037,-0.00507839563851631,-0.0140592773652161,0.00259542948833702,-0.00510119576683066,0.0194104523215852
"2341",-0.00537832281293393,-0.00711474917959598,0,-0.00997148543070703,-0.0059478190975879,-0.00164062816345445,-0.0169821173320315,-0.0112967384234534,0.00378244091970714,-0.0042313265506686
"2342",0,-0.00222379237034187,0.00742597444700399,-0.00604329598200903,-0.00256435682081391,-0.00109560241256357,0.0106815489538958,-0.000714038881167167,-0.0128119161415494,-0.00424916097384553
"2343",-0.00172288202890436,-0.00421020667522631,-0.00655206961672616,-0.00636934991155325,-0.00412891296646711,-0.00109672461534938,0.00626328047292346,0.00905204229746825,0.00288407840261318,-0.000711300967053075
"2344",0.00148603012224835,0.00547116223619093,-0.00412199862600782,0.0107807607123263,-0.00453748862172587,-0.00210459874244306,0.00363089869606004,0.00779033690939346,0.00397525152731326,0.0128112856578488
"2345",0.00205830539274499,0.00469967573404562,-0.000827780680755619,0.0060537812664101,0.00998051660180854,0.00550161017098438,-0.00025875802944153,-0.00163990113413781,0.00286439771350633,0.00913564938547906
"2346",-0.00907583290519953,-0.0051699404422435,-0.0455675120555246,-0.0103153011718328,0.00412370347577573,0.00346541693736979,-0.00232596455267087,-0.0063351757662331,0.0189012095186389,0.00557102644813079
"2347",-0.00539887568168962,-0.00247468104402426,-0.00868057471620687,-0.00434264887098101,0.00255727244989479,-0.000363386360729412,-0.00829025884437673,0.00023645442817255,0.0194575066414584,0.00969530142169384
"2348",0.00794853497621228,0.00744234774756514,0.0183886528952018,-0.00261716483400543,-0.0100680721336752,-0.00290464061339413,0.0133229122126579,0.00873419075114601,-0.00331584305190713,-0.0137173754198485
"2349",-0.00870320174915118,-0.0201918128053595,-0.00945814345492291,-0.0282798593464293,0.0125958648946589,0.00593499193257152,-0.00219140152119524,-0.0109991242697192,-0.00227198153638397,-0.015299103572847
"2350",-0.00557826373064896,-0.0130686325348767,-0.00868057471620687,-0.0162017029100971,0.00548530568007832,0.00181578624206158,0.0134352401666153,-0.00567864353746528,-0.00609954461694495,0.000706277775116781
"2351",-0.000194902590217705,-0.00483861431907673,0.00525396160887981,-0.000304784472448305,0.00668513284225103,0.00271770056899201,0.00382395096337684,-0.000238373929529856,-0.00114556092910212,-0.00988003858289233
"2352",0.00365895934412208,0.00307066430206415,0.00522661933813184,0.00152529254813927,-0.00427401035294084,-0.0023490946536161,0.00977798284313858,0.00166622650928949,0.0090931432784469,0.00641481120450282
"2353",0.000826372111286222,-0.00127541770984008,-0.00086670262411237,-0.0127931855408411,0.00314268773126347,0.00190174480348659,0.00804828598092966,0.000713007525933396,-0.0205390323104401,-0.0219545936385844
"2354",0.0124339052174498,0.0102170996479674,0.0251518244286431,0.0191296930834226,0.0000760136631745567,-0.000180814469473711,0.00187113741401079,0.0121110849005437,0.00273519266083389,0.0246197266652655
"2355",-0.00935478642048415,-0.00581554890305491,-0.0186126483986272,-0.00242192382122397,0.0056545993287489,0.00153701943418816,-0.017805978568139,-0.0114968047683649,0.0094230448977588,0.0233216012391908
"2356",0.000290484771514166,-0.00279750069685325,0.00775860598508404,-0.00273127507829951,-0.0045588493913431,-0.00270833873745879,0.00494392008089917,-0.00617157423183801,-0.00786111182784688,0.0013812676985363
"2357",-0.00871425209826016,-0.0102013207126169,-0.0136868143101708,-0.0179550146983596,0.00969405937906442,0.0038021814621394,-0.00807367169925177,-0.0100306934358491,0.00453941054673446,-0.00137936242976755
"2358",0.00986535381762232,0.0123679284713922,0.0138767427108846,0.0120855268553048,-0.00861820418161163,-0.00360718038588037,0.00788512215667492,0.0123039241622547,0.000739495528218725,0.0110497861959944
"2359",-0.00933363908745843,-0.00865352375934048,-0.00684354570335721,-0.00459289258817952,0.00167776124948649,-0.00135753201837907,-0.0151418888582154,-0.00166830573304921,0.00344825935677506,0.00751355819875688
"2360",0.000292829873747458,0.00333734026025723,0.000861384318629588,-0.00984315724225482,-0.0142356264969975,-0.00806619333098468,-0.013965365915302,-0.00405827147507887,-0.0173457943270676,-0.00745752564579838
"2361",-0.0034651188567445,-0.00614115361257372,-0.00688440041865046,-0.00931956492484953,0.00432436720126916,0.00100501620788407,-0.010784721854725,-0.0105466161037607,-0.001915029174272,-0.00273227328300718
"2362",0.00631756763381697,0.00823885924751466,0.00693212393557463,0.0100344910851486,0.000769194748641233,0.000639414261673465,0.00801257990788851,0.00436044240428179,-0.00133481268036673,0.00410953283883031
"2363",-0.00136259130669802,-0.00306430384067746,-0.00430270380068842,-0.00186269401171069,0.00222788553319697,0.000638322720174278,0.000912223270713719,-0.00024092696299749,-0.0028401637527371,-0.00545702180239194
"2364",0.0129622158996758,0.0197235354601388,0.00777851202617685,0.0102641921141275,-0.00444605286460409,-0.00164108617930014,0.0119774472678933,0.0125451314959486,-0.0173410400266136,0
"2365",0.00678317447171484,0.0113034717593437,0.00686106108225149,0.0120074573517086,-0.00377362810116122,-0.000456422758025155,0.00154365562352554,0.00309693910580511,-0.00272804767106449,0.0116597902841575
"2366",0.000286626103783716,0.00372585200904596,-0.000851593021816477,0.0066929858126803,0.00517904533991809,0.00310592858963243,0.000642645354540505,0,-0.00341939639033861,-0.000677887099525876
"2367",0.00429922806637162,-0.00247468104402426,-0.00255746282970903,-0.000302087691086195,-0.00146097616788321,-0.00191244232595789,0.00436434790857843,-0.00118732307175851,-0.00823467990676474,0.00407050060119052
"2368",-0.00190252378453137,-0.00843469848100453,0.00769208371995633,0.00120908149523014,0.0023872910074052,0.00118612786023498,0.000128049783268969,-0.00784764488632861,0.00380552662673783,-0.00608106773660633
"2369",0.00204943704995797,-0.00125084756221738,-0.000848233319661662,-0.000603794093500198,0.00405726179868271,-0.000337773119386875,0.000639016316247298,0.00143806735560914,-0.00103391351083759,0.0101970756409457
"2370",0.00304352909292116,0.00300605090337558,-0.00848882393872685,0.0081569918926323,0.00720736270672262,0.00310429520011057,0.00536370884213389,-0.000957271842675134,-0.00232882521426903,0.00201895364593252
"2371",-0.00298701043397021,0.00549441978372589,0.00428087761804496,0.0152832956465059,0.0142357470172463,0.0092836607972322,0.00304894496857888,0.0162911698911015,0.0277513534667821,0.00671589392978178
"2372",0.00508853839290424,0.00322906041699733,0.0102300814451564,0.0106257272858286,-0.00743094273768996,-0.00261514112256966,-0.00620589585206932,0.00660073605977596,0.000336482175382402,0.0120079785873621
"2373",0.00156113492199639,0.00693244221995948,0.00675105185348812,0.00905365801531155,0.00242026677001794,0.00144661655552514,0.00611709423755702,0.00491793489216885,-0.00084088464246368,0.00988800541244195
"2374",0.00325967638207092,0.00221296891594758,0.00586756949568001,0.00723591879669216,0.00535604874482298,0.00117368359176839,0.00531977248310112,0.004660744069795,0.0148123379902374,0.0169711811449773
"2375",-0.0013654070810919,-0.0144750428150842,-0.0116666839127181,-0.0114940139286668,0.00645269378982105,0.001533038020191,0.00151199519973089,-0.00347915851615022,0.00555646034903878,-0.00192551936769392
"2376",-0.00947751517750905,-0.0343539999690158,-0.0177066259723069,-0.0252907850451543,0.00484621119630391,0.00351160798791872,-0.00490633401123364,-0.0188549853331591,0.00404122061855672,-0.0122186152959649
"2377",-0.00771175834090232,-0.0152100600430124,-0.0180258947907345,-0.0140172462395275,0.0044517458304687,0.00197399443712887,-0.000758570707031225,-0.00972688991122073,0.00739281267279135,0
"2378",-0.00196702699254281,-0.0185863808500795,-0.00437042777332419,-0.00332744251144357,-0.000738390504353648,-0.000268490651451736,-0.00544024716859692,-0.012937571151816,0.00105999674706458,-0.00651046168649383
"2379",-0.00139382571114754,0.00533461184685269,0.00965762569610695,0.0106223297153125,0.00384381509603715,0.00304532232378718,0.00915918769148028,0.00339816192394604,0.00741225887624641,-0.00524239253493219
"2380",0.00298412118463021,0.00716385013798759,-0.00434781230939274,-0.00360377552538149,0.00485952408727286,0.00107163779917641,0.00504206303262711,-0.00072554770492872,-0.0105110203751617,-0.0171278363614298
"2381",-0.0037240645458092,0.0150156167025663,-0.00174667689587027,0.00271250786513288,-0.00622948120109978,-0.00338957606290369,-0.0015050509835417,0.00383304244146876,0.012828893924552,0.0234584695446547
"2382",0.00644012023601248,0.0254348958611432,0.0227470028183387,0.0177336503448142,-0.0106916082518758,-0.0042966422643419,0.00188440283725599,0.0248051179501381,-0.0059701332626898,0.00916831322138223
"2383",0.00283856212356737,0.0102056450090249,0.00684361497749286,0.0076788498421354,-0.00462150475058498,-0.00224754150219586,0.00411157061232115,0.00783102261061552,-0.0192354761726765,-0.00778717815876662
"2384",-0.00163099715503723,0.00205132077083792,-0.00924832951960608,0.0025400792567627,0.00164732208670415,0.00198240035910313,-0.00050381170118341,-0.00306120404121468,0.000496573998562511,-0.0058862543246091
"2385",0.0130223283557689,0.0307063090577189,0.022472086717279,0.0241602357864423,-0.0114381183292682,-0.0047663445297027,0.00668071414740101,0.0174776974424009,-0.00653433405236836,0.00789483252926959
"2386",-0.0359090003835504,-0.109483700115075,-0.0414201641585411,-0.0607018542052709,0.0268468925526111,0.0138238596572495,-0.0121462046353654,-0.0733519494909414,0.0490383727496597,-0.0202349783501855
"2387",-0.0179099691521628,-0.0231392473699517,-0.00529095355631959,-0.0128636964045364,0.0249674918148293,0.00864488739111402,-0.00190124088313059,-0.0230460047360466,0.00539682539682551,-0.00199870871444952
"2388",0.01803627792122,0.032248954905133,0.0150707500970522,0.0294755788899366,0.00208333470574096,-0.000176462081636797,0.0217166567973857,0.035897577330821,-0.0107357120303128,0.0160213488817786
"2389",0.0170273292187313,0.0221177952019642,0.0131006609907662,0.0253166683576513,-0.00767244859947325,-0.00406524230610705,0.0128032136520289,0.0175741186349212,0.00414934567507186,0.014454602712451
"2390",0.0136455539533682,0.0221801886150179,-0.0086209046183463,0.00999402204362987,0.00368509095881464,0.00221812681459399,0.0111683715372597,0.00827051413379998,0.00500639717121421,-0.00582893627845582
"2391",0.00210069387860212,0,-0.0017389738894239,0.00960403130124243,0.0138847604571726,0.00264209567918572,-0.000728305146817987,0.000482582469987003,0.0153396298304764,0.0123778149562057
"2392",-0.00719345686049266,-0.028314261728461,0,-0.0213316639217349,0.0125202613214372,0.00548238515082433,0.00765215124560203,-0.021702305375958,0.00825478519570799,-0.0283139731648793
"2393",0.00599795338961995,-0.00408520311733973,0,-0.00265104474091871,0.00161578973147503,0.000175679361406056,-0.00361594702129509,-0.0014789891805379,0.00587004706982275,0.0039734554960511
"2394",-0.000620129062908426,-0.00519543895277008,0.000871001593740983,-0.00265796259251572,-0.0000695042218306074,-0.00131861480753137,-0.00883150928188869,-0.00271540505645995,-0.00376250491476637,-0.0283641363814513
"2395",0.0148904159289687,0.0156680236579472,0.00696248500400842,0.0216169415560172,0.00736583265832014,0.00193695185558496,0.0147686604018986,0.01683156070865,0.0060120161086783,0.0101833702572474
"2396",0.00352703078593208,0.0135320696091568,0.02420056275878,0.00956518442475285,-0.0087745345002409,-0.00527292469032181,0.00721668243660512,0.0131452083361203,-0.00942392707864148,-0.00403234117737061
"2397",0.00726319525342056,0.0149528646416253,0.00590722872717131,0.0140685031086385,-0.0164398124831819,-0.00591808915984482,0.0011940840971032,0.00937006929659256,-0.0165518687900309,0.0188934773809963
"2398",-0.000139545589486922,0.000263350026818321,-0.00167790339390939,-0.00169893347202854,0.0117855775061582,0.00257679742937555,0.00417486273691603,-0.0021420833352106,0.00920176941876893,-0.0125828817108378
"2399",0.0055833854320182,0.0105205945081899,0.00168072348555004,0.0144640873147972,-0.0145431367467584,-0.00416589093327024,-0.00736463554179856,0.00620223766322048,-0.00771512582601408,0.00402422820351811
"2400",-0.00134175024871386,-0.00598649872352108,-0.00335578431900785,-0.00223665568237918,-0.00859592342768367,-0.00382734027783649,0.000837883824804209,-0.0111425923787148,-0.00384831534048036,-0.00267204288248979
"2401",0.00268733223598772,0.0023567334819492,0.00252547609119991,0.0089658834103834,-0.000939759270160212,-0.000267951185030646,0.00251079892510364,0.00311691976122308,0.00157682912572787,-0.00468862042717499
"2402",-0.0010165942272683,-0.0094044784577364,-0.00671711296415034,-0.0102748003807641,0.00564166653263043,0.00268131305955022,0.00453179585258257,-0.00286809910742336,0.00133814545546174,-0.00605644537272443
"2403",0.00416299335503201,0.00870254205509102,0.00845302495884948,0.00505070276522557,-0.00546597450929998,-0.00205019675562312,-0.000237419268918737,0.0105461949476811,-0.0143070514449103,-0.00677045791683872
"2404",-0.00377708471671867,-0.00235280367886059,-0.00754402283288347,-0.00307105171507105,0.00202493891185385,0.0022328340229989,0.00142501903472536,-0.00189741970055002,0.0152325067009531,-0.00545330161916657
"2405",0.00448501996525907,0.00183430653153027,0.00168924058233721,0.00728084946155949,0.00173193957522622,-0.000802229240375429,0.00830087845393734,-0.000712850131790344,-0.00746272566859252,-0.0020562452815841
"2406",-0.00271586314845407,-0.000261572324966264,-0.00337267080913661,-0.0100083375265605,-0.000720328278355109,-0.000802805777773585,-0.000940987224878009,0.00356722784420715,-0.0069647567386586,-0.0109890024443174
"2407",0.000461750816527218,0.00340150475346124,0.000846038046968589,0.00786293382861913,0.00158616185151339,0.000624692625094125,-0.00459082514577747,0.00545016871064874,0.00422410931518202,-0.00416660978580086
"2408",-0.00106138697810654,0.00651864190797768,0.0016904872650858,0.00334341718086639,0.0124531598470792,0.00428226702176815,-0.00709579480585754,-0.00023577968394406,0.0161111031746033,-0.00976298245846985
"2409",0.00115461152492746,-0.000518043553628167,0,0.000277699763811201,-0.00184920074104422,0.00053306820047605,0.00738459110991196,0.00495072553354281,-0.00288990863774041,-0.00281693550467965
"2410",0.00161462495718689,0.00959054848212526,0.0177215957753563,0.00527501240322503,0.00833430277101099,0.00381748622955635,0.00969503215421263,0.00680237718361321,0.010339902543008,0.00847467913859545
"2411",-0.000829050387929131,-0.0107833577641967,0.00331673938373123,-0.00193310097479915,-0.0108416948479747,-0.0034718882018776,0.00351263386654255,-0.00582467401828357,0.00186079242861803,-0.0175070513551416
"2412",-0.00640724189156772,-0.00259515515925213,-0.0123965732064955,-0.0071942202830394,-0.0103027195050125,-0.00239949780940729,-0.0151687778652748,-0.000937202363453293,0.00812570029309945,-0.0014254239409307
"2413",0.0029226474867694,-0.00416352149604282,-0.00502102776277891,0.00334447021687301,0.000578205727788994,0.000534542779285108,-0.00426541833718386,-0.00821023437279433,-0.00475942259125139,0.0164167665089441
"2414",0.00106403022317014,0.00418092888332189,0.0142977245616296,0.00555547609743523,0.0075140323519518,0.00240391687275876,-0.00238018019955932,0.0070952739102188,0.00169688399677059,0.0042135701416901
"2415",0.00817900368429014,0.00338283042432996,0.00331673938373123,0.0116021714859131,-0.0103978394798372,-0.00621768184189064,0.00131203929607793,0.00234860227799483,-0.0178639569517192,0.00419567454347969
"2416",-0.000595917816195946,0.00103719060932805,0.00413216893426793,0.00710004127536101,0.00188370784034797,-0.000536455434623107,0.00095320352387418,0.0023429769322274,-0.000862414719033699,0.00557102644813079
"2417",0.000596273145986981,0.00958537819401051,0.00905363056610198,0.0067787485865034,0.00983638623859684,0.00357707490002612,0.00368899812756829,-0.00233750022312551,0.00408032793345359,-0.00277004539170966
"2418",-0.00247513700296464,0.00384930956030138,0.00326254512992641,0.000269293707182428,0.00386743081595409,0.00267351577506103,-0.0013042608763576,0.00421740129612913,0.00468895752335863,-0.0118056088131202
"2419",0.00464079721539901,0.0079242073778456,0.00731717614890748,0.0129239690642922,-0.008917562073118,-0.00479908204048995,-0.00949766501719196,0.000233261940580931,-0.0069228376932613,0.0154603742383221
"2420",-0.000869074720424745,-0.000760665802181815,-0.00484274031442211,-0.00372129670026689,0.00842254790283858,0.00357196331690424,0.00275660609776329,-0.00186587347886424,-0.00211479599145925,0.00761242387006322
"2421",0.00288387045590754,0.00203029721168901,0.00567717665507406,0.0104054271792982,-0.00942380329896786,-0.00293620010036821,-0.000717138370098347,0.00397276300770999,0.00345364201799625,0.0164835036664763
"2422",-0.00515756400749456,0.000506496498135833,-0.008870925101226,-0.00448888281796089,-0.00266595453145924,-0.00169609989882324,-0.0117224192446284,-0.00256054658052618,0.00492807430938913,0.00810813667656118
"2423",0.00188104615263462,-0.00151888943753087,0.00813681354877005,-0.00636617068639589,0.00599711161644945,0.00160915222071933,0.00290487215873747,-0.000233468686682725,0.000233509767000095,0.0040214617765566
"2424",0.00224384941120892,0.00760690347096538,-0.00484274031442211,0.00934332701557183,0.0015805438024652,0.00178528125593269,-0.00289645831761165,0.00373496968586018,0.00474708949416347,0.0126835420999869
"2425",-0.00146207899737805,-0.00830420708509572,-0.00243306640002883,-0.00555401009020562,-0.00523484891857706,-0.00338580365398078,-0.00726220143576628,-0.00697674362126943,-0.00882968004934037,-0.00329593395865624
"2426",-0.0000458537218986921,0,0.00569102329262949,-0.0132978562138598,0.00843457308887618,0.00223495349463643,0.0051207810445002,-0.00210768231034719,-0.00148473859900955,-0.00925926871340432
"2427",0.00201346905571276,0.00456729912620224,0.000808442898791784,-0.00404299528081498,0.00107247363691143,-0.0000893398780495991,0.00218336523285045,0.00657112445725039,-0.000156495540432733,0.00400528569093561
"2428",-0.0051147754056402,-0.0030309849899488,-0.00080778984682639,0.00270614369873079,-0.00235695514083956,-0.000356639647211887,-0.00484132268904081,-0.00373049349893628,-0.0111146366450433,-0.0119681274213354
"2429",-0.000688663949635848,-0.00430711429775388,-0.00485037592410753,0.000809802234422952,-0.00379345666479725,-0.00160606805685548,0.00364849073284912,0.000468340348255714,-0.000870611077112948,0.00403776877017403
"2430",-0.00188328799839022,-0.00534349163512327,-0.00731114476961736,-0.00863013627701525,-0.00582057315059359,-0.00384357199414642,-0.00933107528352606,-0.0112283417270046,-0.00142596843636289,-0.00335122964418233
"2431",0.00492435769681809,0.00460468817148918,0.00327340008305321,0.00761695010879282,0.0133712795033252,0.00412770831355025,0.00941896434895906,0.000709893042637466,0.00198333989726285,-0.00403491472006745
"2432",-0.0016487543009569,-0.00152801198859398,0,-0.00269971636897859,-0.00385157863626107,-0.0000896443286677595,-0.0016964442456151,-0.00520102695448466,-0.0100554550263946,-0.00945308182100768
"2433",-0.00284391361274627,-0.0017850726716897,0.00163119610503504,-0.0110989247559506,0.00143177606624878,-0.00116186955220676,0.00194241562343334,-0.00166378228105213,-0.00199952013116467,-0.0190865205881448
"2434",0.0000458687166424721,0.00562085444556404,0.00732898452683428,0.00766490638040529,0.00110329170342283,0.00156819417921983,-0.00169635556832459,0.00928370757932218,0.00408720952145547,-0.0111189659261556
"2435",0.00450815976828167,0.0149898435735749,0.00727559636331265,0.0162998031966899,-0.0081564423392273,-0.00259436965447957,0.00800958279877761,0.00117954799120024,0.0102162901251792,0.0112439874393682
"2436",0.00302233913994199,0.00550669447821561,0.00561803090342594,0.0213847020608149,0.00728558533300361,0.00466379854932564,0.00710334317952444,0.014840723231877,0.0169076953464486,0.00694917489634173
"2437",-0.0000912743233583146,-0.0002488566208253,0.00478863221504811,-0.00314064274289505,-0.000716271691657111,0.000535494709519302,0.00573833304918026,-0.00580301011378648,-0.00341856092044179,0.00897172432975935
"2438",-0.00228304274261504,0,-0.00476581050135061,-0.00262515194151935,-0.0125407044727976,-0.00490716214843756,-0.0114109645315328,-0.00256822668346912,-0.00530137973645028,0.0177838964431223
"2439",-0.0239348519871588,-0.0209162033507168,-0.0159616656343274,-0.0336933620639602,-0.0164745437401388,-0.00475193355303272,-0.0397980288484594,-0.0255150099050973,-0.00658355691146817,-0.0154570542315235
"2440",0.0143471758048095,0.00890115683145987,0.00811024305510299,0.00681037926714034,0.00051646041363318,0.000900838191176812,0.0121463062102167,0.0048039547903731,-0.001262358974359,0
"2441",-0.014375454608089,-0.0199140595412522,-0.0176990303820017,-0.025162487631838,-0.0113578844111493,-0.00369047657663013,-0.0243723186606559,-0.0207983925238253,-0.00663556384028952,-0.0129693172763443
"2442",-0.000375012959172083,-0.000514541814449876,-0.00655200854611149,0.00305312250284273,0.00149241282377255,0.00225901234069936,0.00304349294918138,-0.00170886212097188,0.00341948310139162,-0.00760708883651384
"2443",0.00999268173106649,0.00797722549937951,0.00494645400501681,0.0171553879983641,-0.00432104359991736,0.000270023104559369,0.0045513360331928,0.00611396854151036,-0.00641937708036144,0.00487798195622902
"2444",-0.00386538817642135,-0.0178707462713303,-0.00820356298098124,-0.0068007592853726,0.00807998132619381,0.00108125930159764,-0.0010070654271831,-0.0110591936192251,-0.00247272068741999,0.00138694364428016
"2445",0.00018752229446628,0.0077982435677395,0.00330859824608165,0.00794300248918178,-0.00326574804722302,-0.00171025000329983,0.00944813913912701,0.00793480518959688,0.002079018104574,-0.00069244007257252
"2446",0.0000469476939330971,0.00206340402114891,0.0140148352551683,0.00054332822493941,0.003499785965835,0.0015331028026484,-0.00162215143170052,0.00442791852846347,0.000957564634535668,0.00346495601403118
"2447",0.0112452539422838,0.0128701855340903,0.0292683344265299,0.027974222855792,0.0080873112493276,0.00162057418125272,0.0114998793302121,0.00857201449566247,0.0145886078668909,0.0124309117376125
"2448",0.00630152873705425,0.0116900261525561,0.0126381282793091,0.00713316595775293,0.00794871890857207,0.00296627474019595,0.0194020693889037,0.0114133438810065,0.00235721699592717,0.00545709200812983
"2449",-0.00547922383696808,-0.00753586638782311,-0.0140405093775716,-0.0128540173898103,-0.000949252979055237,0.000448043945477705,0.00254580220156031,-0.00408155035660684,0.000627122364192267,-0.0115332945108013
"2450",-0.00810221755551965,-0.0111364616466029,-0.00870257414079834,-0.0146159487240335,0.00635824978509714,0.00286657789122713,0.00117051016680159,0,-0.000783384241545115,0.00686346568920571
"2451",0.00620785512977196,0.00076781717240082,0.0111732899187951,0.0142933708550341,0.0073358214506094,0.00169695744688703,-0.00779532286506435,0.00771450597455203,-0.0072912581585749,-0.00954336553088786
"2452",0.00496362088972901,0.0112533241518136,-0.00157864334840474,0.00904029250864702,-0.00216307699197038,-0.000445720074611633,0.00552413304463339,0.00334928751024943,-0.00315907432098228,0.0233998982825621
"2453",-0.00904724152055314,-0.0144160732380617,-0.00711464035578446,-0.0173914733173268,0.00252898761709019,0.000624450001357246,-0.010743544178422,-0.0164520161740668,-0.00118840911750584,0.00605251050862865
"2454",0.0075461514612456,0.0105211070012206,-0.00159214939101582,0.00429076800783457,-0.00893685127271293,-0.00249649134425123,-0.00481277019859683,0.0111513704686619,-0.00341081145395405,0.00334226902923129
"2455",-0.0024042581755922,-0.00152351754695101,-0.00318978254657198,0.00694247907372958,-0.00330039494478795,-0.0023268145198273,-0.0181051665440006,-0.00455522565842004,-0.00254695162804008,0.0086608425336514
"2456",-0.00509763139844599,0.00152584219430785,-0.00560022322729936,-0.0111375925467742,-0.0116950765089998,-0.00457538685139569,-0.0143976528414501,-0.0139690513441701,-0.0347111315033514,-0.0026419718257199
"2457",0.00442529062542074,0.00253925247328035,0.00643619517625171,0.0144811628482999,-0.00465941141594561,-0.00225301908295805,-0.019349129166241,-0.0134345125903319,-0.0015706538681437,0.00596018324407677
"2458",0.000695382494254604,-0.00607897350945741,-0.00479626590524385,0.000793105221192469,-0.00557303836302969,-0.00207744642972663,0.00169881784235604,-0.0118839988847488,-0.00927301713258011,0.0019750244006882
"2459",-0.00342915040964864,-0.00764522018703007,0,-0.00449041318998877,0.000672888467173616,0.00144824166514934,-0.00143519981907447,-0.00876974562582644,0.000668510758197849,-0.00262808499404299
"2460",0.00520821010400629,0.0023114275866758,0.00321292779591587,0.0108782969133014,-0.00589904286097997,-0.00262101597332898,0.00587857791867563,0,0.00350764996672215,0.011198928205062
"2461",-0.0126295093332506,-0.0148605705457645,-0.00880708817996445,-0.0230973211429709,-0.00225368067832366,-0.000272059861371798,-0.00999987643751077,-0.0171890930083848,-0.00507657273380246,-0.00586324608441957
"2462",0.00131191258290819,-0.00286065894592202,-0.0016155580597087,-0.00188041025704744,0.0009788864456719,0,0.0135116496657475,-0.00154312200135476,0.00158925131938314,-0.00720842462624149
"2463",-0.00327544893333453,-0.00443423246518604,-0.00161808563522059,-0.00888316999272043,0.00376032963246109,0.00208493712893354,0.00556584256561488,0.0108190816621758,0.00242192253920037,0.00660070625287879
"2464",0.000516486853260334,0.00104813832683259,0,0.00162972170593889,-0.0140115179202065,-0.00307527852258593,-0.00334678624658402,-0.002803129815937,-0.00558192123287449,0.000655728765314612
"2465",-0.00347225859238398,-0.00366427875590125,0.000810495116301935,-0.00108456546244518,0.00638343603554681,0.0021775714936636,0.00129138819779206,-0.0053668002414492,0.00268095674697588,0.00131066557908799
"2466",0.00626229902758069,0.0123460094742609,0.00566780858346672,0.0176438348927965,0.0032468651112445,0.00199159844313335,0.00683595993411767,0.0125899805581686,0.00618313836898388,0.00196339129656375
"2467",0.00266711763207628,0.0015566076270046,0.00322060243631861,0.00613486132518393,0.000827981504498254,0.000451940352519387,0.00422793864640814,0.00558223987559692,0.00572997019980015,0.00653165629159558
"2468",-0.00186658397663264,0.000259324726260779,0.00882838033762257,-0.0029161285240108,0.00105329619016414,-0.000903316678711907,-0.00382731995899988,0.002523806656761,-0.00305509864540421,-0.00908501892228064
"2469",0.000467460587354029,-0.00259020966627788,0,-0.000265856832991962,0.00150244303102287,0.00108508670631502,-0.00128060620353487,-0.00226576314927696,0.000745436487418205,0.00392921932243606
"2470",0.00425277943225555,-0.00129835245883569,0.00159113829062152,0.00425527569208528,-0.00435122284000133,-0.00135472036645645,0.00269275228358623,0.00227090849004918,-0.00223457746859923,0.000652373967855002
"2471",-0.00335071645579399,-0.00259999386683263,0.000794209566832071,0.00105949182064458,0.00263739905000859,-0.00018100237923091,-0.00191814100824861,0.00125792861587293,0.0075481338345742,-0.00456323801298775
"2472",-0.00200765921192603,-0.00547443199864739,-0.00158724362195761,-0.0105820887605579,-0.00676339166438933,-0.0021705604458151,-0.0116591212208582,-0.0103067784156486,-0.00559809001730394,-0.00654883367309145
"2473",-0.00266674337554251,0.00183478734145925,0.00158976696944024,-0.00855617861939462,-0.0108937490772314,-0.00344397598656931,-0.0229454217814723,-0.0111755960905677,0.00182135109014525,0.0059327489710721
"2474",-0.00295534525543006,-0.00130832037149431,0.00158743492783686,-0.00404538189595982,-0.00221815180134666,0.000181840344236406,0.00199016363161086,-0.00616515704754228,0.00471035443830492,-0.00655305811402018
"2475",0.0000470636459284357,-0.00104781737586512,0.000792321539675234,0.00568644435178456,0.00613253649513879,0.000818412030803906,0.0148305226907144,0.00749557953344882,0.00296101327585108,-0.0131925678921104
"2476",-0.0072453567930485,-0.00445844985851074,-0.00395883181348788,-0.00807748800811314,0.0000762285298239185,0.0000363806739398509,-0.0220509713326773,-0.00384828944830296,0.00647860412533041,0.00467914912177814
"2477",-0.00601875842768285,-0.0071127742151873,-0.00635921690776942,-0.0119434693491463,0.00435123626292033,0.00300251036118837,-0.0128086407947137,0.000772704509771183,0.00741461727170334,-0.011976089318696
"2478",-0.0045771340501769,-0.00212273716020739,0.00239980488394775,-0.00274739304092442,-0.00767630444215461,-0.000635133025918777,-0.00581170117393037,0.00257318242977034,0.0053381106869792,-0.00336702670285538
"2479",-0.00110180848063168,-0.00904006912342559,-0.0119712171633061,-0.0101928335166621,0.0089606164394469,0.00308603155217746,0.0053017400543891,-0.00769986731696304,0.000724022508671984,-0.00675673420271494
"2480",0.0220572808431472,0.0160986553396589,0.00706776634024786,0.0361814038443713,-0.00850156155047044,-0.0041621482775267,0.0163625296839589,0.00931168565843099,-0.0180078544738954,0.00408164694177549
"2481",0.00450382739826138,0.00316876600723082,-0.00120299837032378,0.00644642232775872,-0.00405751351925654,-0.00354413596169101,0.00612025744335609,0.00256283036433347,-0.0041752189246792,-0.00135499503103398
"2482",0.0106021294558571,0.0050013598044274,-0.00843207758086062,-0.0325593901771768,-0.0424322276445011,-0.0152288451346184,-0.0185134061317622,-0.00434571408479856,-0.000657686621651554,0.00474898719275374
"2483",0.00249559645766051,-0.00366669197625935,0.000809894341520012,-0.0284137299956269,-0.0147708382573254,-0.00601920172939652,-0.0181893379109982,-0.0269576171011647,-0.0148897501627139,-0.00810266141648341
"2484",-0.00230515461053449,-0.00972669124476577,0.0014161789877547,-0.0190233424833495,-0.00562179881296132,-0.00204949237592789,0.00535211475487074,-0.00765178633065577,-0.0221294530271399,-0.0190606052729353
"2485",0.000785668308206366,-0.0082294639021131,0.00121216344814701,-0.00723583468081312,-0.00598186903088249,-0.00578774509837887,0.0169258376958097,-0.0124964425828747,-0.0084542870786386,-0.00208185917709702
"2486",0.007802740926796,0.00588877768782137,0.0016141458945611,0.0201165827023355,0.00494599811994156,0,-0.00362412495320241,0.00700049925425428,0.00869866498407834,0.0222531114282418
"2487",-0.00187850640382281,-0.0119743766074448,-0.00483474178748255,-0.00828796139002197,0.00902316398436542,0.000939018544820591,-0.00215560401548665,-0.0131015898839957,-0.00298843913110214,-0.0122448708106266
"2488",0.00514086233146238,0.00457852646044565,0.0149796855020301,0.00144091725268214,-0.0147145295793185,-0.004409148885269,-0.00823535392605423,0.0149010734736781,-0.00513829763993223,0.00206601655464245
"2489",-0.00223761378167697,-0.0109921559117417,-0.0149581473269729,-0.0046045519266823,-0.00288762058252534,-0.00442813822904531,0.00299478106341566,-0.00854238461867152,-0.00878020158010162,0.0082475228783081
"2490",0.00755156329639561,0.00975895748754874,0.00809883496076425,0.00982961992136322,0.00248231261471332,0.00085161211165663,0.000135758240104256,0.00215403997030261,0.00373425959645224,0.0279482321863713
"2491",0.00195327636830367,0.00107366625348648,0.00241009895819722,0.0151731523730827,-0.000330012126703472,0.000945606906831431,0.017098850222196,0.00537326440100738,-0.000346089282815432,-0.00132631000327676
"2492",0.000543963030960271,-0.00724054213796321,0,-0.0107161413990955,-0.00388080679167768,-0.0035900722144655,-0.00547034550769787,-0.00213771495799142,-0.0198199842494375,0.00398407763104802
"2493",0.00371544481128305,0.00810389597887262,-0.00841518327070734,0.00484589377406808,0.00149214888818117,-0.000853462761718826,0.00509773572381866,0.0013392416552358,-0.00565120529801322,-0.00727510080633487
"2494",-0.00469483082825939,-0.0112542152799887,0.00868858826800389,0.0039716180544882,0.00736618902352837,0.00455523682992021,0.0034705271296358,0.00748819309840676,0.0105674628312986,0.00333106690960094
"2495",0.00195042629994724,0.00840106957439923,0.00100163042590684,0.00141276217460495,0.00419043011494802,0.00103884885496242,0.00824676451145745,0.00398218601130895,-0.00465734609866397,-0.0199203198141998
"2496",-0.00239921414007349,-0.000805838624679756,-0.00160092359739905,0.00169318146945119,-0.016200374010807,-0.00669984783443944,-0.012532715753431,0.000264400983798874,-0.0134192375762137,0.0304878065787826
"2497",-0.00367545009231041,-0.00134503618354909,-0.00841847092918646,-0.0118309148328575,-0.0105585702866787,-0.00381514426244889,-0.0157649792356636,-0.0129526682818182,-0.00187918568232659,0.0184088928598929
"2498",0.000500750981371034,0.00296268710147096,0.00303205144155472,0.0011400914013544,0.007327480392747,0.00448863940362165,0.0105875364873405,0.00723059504786572,0.00537921816945297,0.00710139187360448
"2499",0.00600882125608093,0.0158430638245239,-0.00120905936088511,0.00825746892857304,-0.00108680530792915,-0.00038042240218128,0.00792513603995504,0.00452012163201365,-0.00535043700151983,0.00512820106818124
"2500",0.00316747206230428,0.00978036152699024,0.00443892282652447,0.00536588255673665,-0.000753599937245775,0.000380567178461577,0.00639628644235168,0.00608814191558205,-0.00098620225043744,-0.00446429040277008
"2501",0.0130807238430899,0.0141363797866028,0.0148655111623044,0.0168536888231263,0.00854414798518555,0.00332779448368004,0.0194652122351822,0.0142065551139581,0.0035897155164677,-0.0076874068323729
"2502",0.00244865398610972,-0.00438824685218864,0.0114804786630931,0.00441999538943461,-0.0117940595847199,-0.003790527062706,0.00506542064499693,-0.000778115506416821,-0.00232497536752252,0.00193683988393856
"2503",0.00604039993959504,0.00518521472299982,0.00293548144375833,-0.00522571469253874,-0.0124388297167225,-0.00513632046008539,-0.000775259401985862,0.000778721441645702,-0.0104866720444563,0.0051545684159735
"2504",-0.001147761789415,-0.00154748838277774,-0.00975609664325361,-0.00663522125818672,0.00187225928223089,0.000190765354217248,0.00620789772801911,-0.00544724489646586,0.00380432964122579,0.00641030081676885
"2505",0.00667399802687285,0.0116247409015393,0.0118225449835323,0.0111328424042636,0.00356775341614157,0.000573635171625897,0,0.00808529674364378,-0.00333877458942422,0.00254773579355727
"2506",-0.00825417637573844,-0.0145556256278959,-0.0153845142794972,-0.0297276063635333,-0.0111730897337152,-0.00831156581922943,-0.0185089254191836,-0.0165586120604729,-0.0146672253870682,-0.00952992615734338
"2507",0.0041172273697796,-0.000259045607986619,0,0.00170230770263879,0.00505046094533745,-0.00279400800169893,-0.00746481003072397,-0.0144700088905011,-0.013691132708056,-0.00128285619031576
"2508",-0.00195600825618303,0.00311044971675867,-0.00870257414079834,-0.00453127843209444,-0.00229989917573503,0.0012559905960825,0.0133264848936367,0.000739237183633668,0.00661456145386863,0.00449589628991709
"2509",0.00217743757968147,-0.00361753847436896,0.00857928893802651,-0.0068279807056757,0.0107566313816632,0.00463171987982203,0.0110677556151657,0,0.00499762133278225,-0.00575452855061109
"2510",0.00385777659096176,0.00363067257208627,0.000989232084672498,0.00343727378441905,-0.00498292642023435,-0.00211311277574466,0.00180290973833319,0.00653393536837599,-0.00736711510699384,0.00450167871434171
"2511",-0.00278276780078268,0.00155037363187249,-0.00533818746800097,-0.00415749748708472,0.00441349434360294,0.00163614696020886,-0.0123055354938719,0.00028229666581292,0.000556610069982311,-0.00576196249489347
"2512",-0.00172753860972663,-0.00179361402379008,-0.00160799478412244,-0.0118876373574829,-0.00178742387645725,-0.000433170997025889,-0.0018476308316886,-0.00395048942982157,-0.00241077426816461,-0.00128774623731354
"2513",0.00146433630248555,0.00286438068497241,0.00181195297544123,0.00586838911402299,0.00203691267676986,0.000962922962444601,0.0026441550718026,0.0048160633792218,0.00316018229055426,0.00193420953618118
"2514",0.00248098158776111,0.00129856471887901,-0.00622995877233168,0.00437592865465586,-0.00321870578155459,-0.00144318069620386,0.00118685516436834,0.00535642285192872,0.00583709811915112,0.015444003425422
"2515",-0.00826447731962432,-0.00622429321553308,-0.00141546440421925,0.00755136599775863,0.00730842887082606,0.0036608374369218,-0.00592689774851707,-0.00701043345287511,0.00276347646948194,0.000633704922959666
"2516",-0.000222895778161925,0.00704618740392826,-0.0101255541522219,0.0164313996990675,0.00354317232679713,0.00307135895736343,0.00993751429890977,0.0104489878211058,0.0131361380384334,0.00126673755373652
"2517",-0.00365490161981896,0.00570098499134475,-0.000409180788950025,-0.00709030516086118,0.00151332558474082,0.00296601894947668,0.00944625673032196,0.008384698326249,-0.00616556345846808,0.0018974420434541
"2518",0.00765001905177431,0.00231893193277855,0.00818670564552981,0.0119966194227066,0.00428133629802541,-0.000476704054778621,0.00402923079358875,0.000831430623377871,0.00784599938102359,-0.0119949157764663
"2519",0.00594936106498567,0.00874015751611323,0.0200972884663349,0.00762066605059641,0.00384472358711729,0.00114501219422025,0.0137217136574637,0.0105234458930408,0.00353037020430547,0.00766769250680732
"2520",-0.000794483424922943,0.00866485157153707,0.00577126854614063,0.0109244012029188,0.0156534455153936,0.00648322831630344,0.00344780507498732,0.0150725587353084,0.0155150729251752,0.00507298460463712
"2521",0.0035776695261498,-0.004295068808707,-0.00158300643534548,-0.00415625563137267,-0.00918162913250953,-0.00454681553667291,-0.00216334766706017,-0.000270026178959326,-0.00737255272033122,-0.00126187729913718
"2522",-0.00330079669700412,-0.00380630714835262,0.000991015904208359,-0.000834738443369454,0.00802583103328791,0.00380627364316855,-0.00663189778472451,-0.00189052973516601,0.00823264429530202,-0.0151611396094232
"2523",0,0,-0.00376180504080792,0.00584784045578712,-0.000656844285984115,-0.000473818666142933,-0.00937224520898661,-0.000540925563579986,0.00426026456483997,-0.00448993064839287
"2524",0.00282608454166078,0.00534895417411962,0.00655816198224479,0.0119049019611941,0.00336761793924012,0.00113788903722534,-0.00427656983438574,-0.00243632116655024,0.00309322133286405,0.0109535241994081
"2525",-0.00251008547511211,0.00177358237679903,-0.00157931764186536,0.00437754930891798,-0.00221014778286566,0.000568262288961563,0.00455520091718475,-0.00407078191786148,0.0036123700440529,0.0146590152638848
"2526",0.00229575357606948,0.0037935973735328,0.00632764025799815,-0.000817229630920235,-0.00475840083618828,-0.00217752143282135,-0.00103637727245365,-0.00108994580529775,0.00263361416438879,-0.00188439640516536
"2527",-0.00352362919261162,-0.000755885495406283,-0.0112006894268618,-0.000545353572565688,0.0104691647107409,0.0050287788790675,0.0067445800762449,0.000272891482451687,0.0143595045474083,-0.000629382790976241
"2528",0.0022098919427791,-0.00378211923034433,-0.000198598898137003,-0.00545554059650999,-0.012808169958276,-0.00708085925607216,0.00167474302375181,0.00054533586911143,-0.00845917148828956,-0.008816065726727
"2529",-0.00370443945592014,-0.00253089205454149,-0.00278278916697983,-0.00301687805214279,-0.00685883285706401,-0.00380292031410123,-0.0104181476613501,-0.00981178831254226,-0.000870601526840709,-0.00317664205244783
"2530",0.0036740471850456,0.00532839808154106,0.00637840770999065,0.00192551683360009,-0.00199702521146206,0.00047693140991556,0.00636869578920884,0.00385364457859128,0.00243971427480294,0.0114722499988849
"2531",-0.00260215095077054,0.00328139348982392,0.00059414709322736,0.0148271198918624,0.0100051246730843,0.00524704012202837,0.00762002115791183,0.00795168198175999,0.00643196854153927,0
"2532",0.00641173080897084,0.00201246643595177,0.00257322039307772,0.00622296041365744,-0.00685187565483791,-0.00379617006936395,0.00230696375213202,0.00108816657928856,-0.00449092318429123,0.00252050941723025
"2533",0.00865548433099028,0.0120510468190036,0.0104640195300318,0.0110244794159362,-0.0125507086006449,-0.00495346691789111,-0.00537112959481267,0.000543376324157796,-0.00824149409841668,-0.00628526933019513
"2534",-0.00104532902583565,-0.00620168702471258,0.00136770105097872,-0.00425533294186742,0.00336699549370501,0.00134019355991422,-0.00102838265916683,-0.00461698237896435,-0.009272200839748,0.00442745156679414
"2535",-0.00156991756901614,-0.000499223310839736,-0.00819516330104819,0.000801324269230408,0.0036074116143987,0.00124315299128974,-0.00939517788551147,-0.00136446474851504,0.00203069041090065,-0.00818635137568224
"2536",-0.00620168443805991,-0.00874139266824481,-0.00275432075917981,-0.00533757738992136,-0.00300945545908016,-0.00028667656525827,-0.00688536691915986,-0.00109272464218724,0.00422947403699836,-0.00571427301828686
"2537",-0.0000879080361245732,0.00377926038127629,-0.00236712809731621,0.00187830433050329,0.00695916899391902,0.00343883037999326,0.00784899963557195,0.00957337020476579,0.0138633147857918,0.00574711359443247
"2538",0.000395656331741101,0.00326305121298831,0.00533901059846764,0.000535483083642152,-0.00618324037378593,-0.00191648861150229,-0.0118119757657743,0.00189641263616291,-0.00302904362538192,0.0107936340731034
"2539",0.000658925853124659,-0.00100072260429585,-0.000393405911207623,0.00428278444442243,-0.000419899277294022,0.000382349575538621,0.0111650477127438,-0.00243358740945254,0.00555554701967576,0
"2540",0.00689292507586292,0.00400692789470303,0.0045257297184369,0.00612984926282567,-0.00041993870045498,0.000763547743473092,0.00675497598482644,0.00542136251197944,0.00250346175771621,-0.000628132135055082
"2541",-0.001787868934498,-0.00947861549086293,-0.00156702599926861,-0.00238408880286523,0.00605068088338445,0.00477074502833719,-0.00335487739760021,-0.00188747146632151,0.0135193321325926,-0.00628526933019513
"2542",0.0000437945892688418,-0.00125912829742159,-0.000588634945132505,-0.00504508206380994,0.00735040078410387,0.00180394459608713,-0.00142396848769366,0.00216111441405342,-0.00203906547253352,-0.00442764686394759
"2543",0.00131046919429667,0.00252140353010999,0.00294455479592526,0.0061381449169704,0.0135984446414505,0.00407576917314612,0.00726047304423805,0.00539084043448312,0.00621490725536278,0.00381195738522355
"2544",0.00593259961752213,0.00402417155075585,-0.00137002769820127,0.00450944536943121,-0.011534477974294,-0.0059472695963152,0.00308928975040756,0.00428961973977526,-0.00761486576504167,0.0050632218761828
"2545",0.00394609065819407,0,0.00705607451126999,0.00924209853590519,-0.000579379185845941,-0.0006646482199405,0.00769903143243811,0.00106770274602863,0.00264299597030426,0.0107053384040592
"2546",0.00544262190377132,0.00450901666272796,0.00389254761451863,0.00313974156893049,-0.00314710563123144,-0.00152045063515105,0.00331088912207567,-0.00293294562619995,-0.00680267868712037,-0.0112149924655612
"2547",0.00399545219807962,0.00074823970716964,-0.00717337899289039,0.00104337045395408,-0.00722681038443673,-0.00361668121522118,-0.00558449687025786,0.000267173501275808,0.00111298798511172,0.00126028713508397
"2548",0.0052201486031882,0.00274100768845043,-0.00097635712399502,0.00807697640483807,-0.00460203642094537,-0.00191024381315852,-0.000893452760813096,0.00187153420193842,0.00444707944924305,0.00125863603933829
"2549",-0.000851154276010901,0.00472169589239302,0.0011728149929886,-0.00361828783326679,0.00546396280500283,0.00401911993084059,0.00472651306633165,0.00080065261034723,0.00536402738264852,-0.00628526933019513
"2550",0.00157630661285846,-0.00321554229902843,-0.000585679204801126,-0.00415057842143496,0.00593579176500669,0.00266926269103585,0.00165312787432104,-0.00106656397274618,-0.0033875507556308,-0.00189763734060744
"2551",0.00595514977644229,0.00124080419383543,0.0084000754083926,0.0109403905354675,-0.00174529763591624,-0.000475316388294456,0.0125665286663676,-0.00240269606376431,0.000594833446634802,-0.00126734462309919
"2552",-0.000888038866522334,0,0.00116244571652979,0.00309203789958512,0.00166528350845585,0.00161696852561599,-0.00250725232729276,0.00240848291618678,0.00135884501061567,-0.00507620312805912
"2553",0.000677071295172915,0.00272617264350217,-0.000967702949906002,0.00025670932937838,0.00299205525868307,0.00265881780106692,0.00427296280120859,0.00453793938462188,0.00873545895223615,0.00318873197427805
"2554",0.00126897325605135,-0.00889775527251324,-0.0021304507809875,-0.0118130768228339,0.0111048170706005,0.00464053940276421,0.00500573381192915,-0.00212582350234125,0.00638973421238043,-0.00190709233946518
"2555",0.00156292023699911,0.00174549755818054,-0.00310556376252358,-0.00311844318660925,-0.00590108005737222,-0.00358208459684939,0.00522968821513659,-0.00399457226108579,-0.00484539694683539,-0.00254780134871879
"2556",-0.00269914877765076,-0.00174245610530355,-0.00253115563076189,-0.00964539991355429,0.00371013230424788,-0.00047302292313256,-0.00396397274001992,0,0.000923438526105436,0.00383143097049166
"2557",0.0139975051101182,0.0117207773941803,0.0117119173032265,0.0155304051588157,-0.0167561060359916,-0.00696660382529646,-0.00310886043968317,0.000801988627725292,-0.00142585755030133,0.00445286527660071
"2558",-0.00629740224836206,-0.00369736636583151,-0.00945394320548387,-0.0176258098019774,-0.00359955875567997,-0.00286350536616264,-0.0041167297451189,-0.0125568220567593,-0.0124306738187582,-0.0158327854283856
"2559",0.00062954582803898,0.00841167462709058,0.000584310198584959,0.00765170057062425,0.00260400123261784,0.000957273576400741,-0.00238018298475573,0.00405860181441997,-0.000595339333299139,0.0051480673719293
"2560",-0.00297793945463776,-0.00515213535330061,-0.00233602022007018,0.000523790782366751,-0.00477571624039419,-0.000191525305466289,-0.0046460125805442,-0.00161680643160456,-0.00672284049488825,-0.00128045807361343
"2561",-0.0029868972995224,-0.005671980904985,-0.00234151065084642,0.00104680732656748,-0.00303076278760894,-0.00143465333663395,-0.00428903425510763,-0.00485843814957099,-0.00805347834087144,-0.00448725015697193
"2562",-0.00185651821385779,-0.00421610396936023,-0.0031292311274409,-0.00941175236556335,-0.00540472082924925,-0.00335213579841132,-0.0153299374194131,-0.00867903284016802,-0.00621869931092334,-0.0225369177448197
"2563",0.00126812056620285,0.00796991541863701,0,-0.00791767435864299,-0.00798084180120184,-0.00278716590448491,-0.0127381388851198,0.000547059808659212,-0.0051277334456411,-0.00856391818071489
"2564",0.00350426482897248,0.00889544814687149,0.00725922847643523,0.0111732558472162,0.00350935182711343,0.00212018340311171,-0.00247622790346769,0.000273729196672345,0.00218397831585593,-0.00930240351013967
"2565",0.000504739138693866,0.00391882153753809,0.00506403547213385,0.0139437318582647,-0.00631155077381262,-0.00250059263465241,0.0015677938637102,0.00191355394184733,0.000174311365286783,-0.00134129435353814
"2566",-0.00382651994140704,-0.00731901709399407,-0.00697645524597157,-0.00570842154139328,0.00480623055830343,0.0010605729410238,-0.000913267590523126,-0.00818579395909336,-0.00540347752141324,-0.00402956400638621
"2567",0.00865358579059583,0.0135169399579249,0.0101481670498955,0.0260959327197492,0.0122152299783973,0.00876443036863739,0.0184099985815678,0.0159560035026385,0.0186645368384717,0.00876603378785168
"2568",-0.00196710702652847,0.0104268200982149,-0.00193202606382603,0.00610372896824396,-0.00506346887830589,-0.00276880511502464,-0.00166668567401851,0.0119145041402662,0.00412905806451613,-0.00133694889041081
"2569",-0.0017562374272041,0.00191973954440638,0.00329084117194922,-0.00176927566760388,0.00627647113399354,0.00268093236474032,0.00423779450164452,0.00263645956555147,0.0022273193979101,0.00334674345417874
"2570",-0.00109681542203477,-0.0019160612059399,0.000192894668396226,0.0116484386071853,0.00429880478375466,0.00238675687398326,-0.000383961595088134,0.000804899647445456,0.00444485861090449,-0.000667102292611355
"2571",-0.0128394499260324,-0.00359979016874357,-0.00771609632218306,-0.0110138156821425,0.00830883022692541,0.00333377847702865,-0.00319783093254167,-0.00750680845812146,0.00876520281226778,-0.00534051833327187
"2572",0.0023530870834958,0,0.00136078823073094,0.00480896217787974,0.00399543808373215,0.00189914927800783,0.000513274599598601,0.00270141160337389,0.00244643999960825,-0.000671062731966487
"2573",-0.0010670807566896,0.00120423853629337,0.00077663936549488,0.000251839029382417,-0.0014093678305489,-0.00104247358399601,0.00743956480991437,0.00404092371710152,-0.00134649497018424,-0.00201488568513231
"2574",-0.00072641250522687,0.00360852980921211,0.00620743053103712,0.00251840807081272,0.00356972378523479,0.000569080669376554,-0.000707016749153633,0.00295139598789529,0.00160110392855994,0.00336476113458128
"2575",-0.0010262383776739,0.00527308875966903,0.000578503243311435,-0.00276322476571544,0.00455017267465085,0.00246503283805,-0.00681727394834086,-0.000534923712668722,0.00563686685481346,-0.00134129435353814
"2576",0.00727687802210375,0.000238488495809541,0.00847779544019156,0.00277088133363956,-0.00667051016781772,-0.00340458565914226,0.00440339027702663,-0.000802960583149548,-0.00409937257675375,0.00604431144893303
"2577",0.000934820556610427,-0.000953463040949565,-0.00133738908816683,0.00175835418719972,0.00596926665145814,0.00284669648060687,0.00438408543783608,0.00267858903233753,0.00243616429405091,0.00934580402420737
"2578",0.00318418996562619,-0.00381783486456488,-0.00554815337152426,-0.00526593863651037,-0.00807679278839935,-0.00283861580299072,0.00295307249536036,-0.00534315731477186,-0.0072069134801489,0.00396826774429404
"2579",-0.00232766575267029,0.00239510298259771,-0.00923438559281509,-0.00705826666242548,0.00290810877819059,0.00199287329580233,0.00473619691383598,0.00456622546126551,0.00211023886122863,0.00197625751826047
"2580",-0.00173913397580927,-0.00382309807414372,0.00504863251140764,0.00558515781685109,0.010086564964215,0.00492246704868937,0.000891808038945285,-0.00106950140172324,0.0053065784593449,-0.00394485458956617
"2581",0.000637420776040676,0.00143922018303022,-0.00347757735351928,0.000505122056369434,-0.00542426459082401,-0.00141548963741456,-0.000891013426009168,0.00214132526797139,0.0022622958066576,0.00990112731437764
"2582",-0.00297275507703854,-0.00670645249734492,-0.00697946726278287,-0.00302816804814077,0.00305771167636015,0.00189024716616371,0.000254973900139399,-0.00160268339233294,0,0.00196069013709699
"2583",0.00281112171262854,0.00337598627855895,-0.00507614832396164,-0.00177170566695772,-0.00148305313407771,-0.000660586684285924,0.00687802270064597,0.00909580465911608,-0.00367833965026731,0.00260929445926572
"2584",-0.0010192833422894,-0.00144230571276049,0.00215862711166093,-0.00177485017907797,-0.00404291310029925,-0.00302051744519238,0.0011386578992767,0,0.00234937909045141,0.00260250376062299
"2585",0.00059511702966053,-0.000962535803794129,-0.00234974271520982,-0.00406391167209352,0.00463919351517639,0.00179904683194376,0.00694955311567247,-0.00397664616298099,0,0.00778704458108392
"2586",-0.00118973964626201,0.00602269663814137,0.00510296508963148,-0.00229542597109578,0.00948306482884687,0.00463118177633781,0.00552147775873935,0.00904986894944892,0.0144818601580603,0.00193185131067319
"2587",-0.00438184913632433,-0.00119742347099827,-0.00331959354262235,0.00485687672108459,0.00547287318652168,0.00310458394125623,-0.00224638363877316,0.00580310799561246,0.00684870852630226,0
"2588",-0.00649492086796255,-0.00695266145958839,-0.00842469988256733,-0.00432464404264055,0.00308716552243493,0.00300172125839926,-0.00200124990374406,-0.00209798827418783,0.00475332744025558,0.00321332361178372
"2589",0.00885988123054671,0.0062771586142194,0.0106696662361043,0.0104753372698998,-0.00307766426343126,-0.00158967352615802,0.0125329636864224,0.0113007444535693,-0.00293637851445971,-0.00576545622459146
"2590",-0.00298421508519175,-0.00527846823858635,-0.00312794567972496,-0.0126424349875188,0.0130797421358055,0.00571300588901824,0.00235195910987462,0.000519789289042949,0.00474478083679286,-0.00386605894290903
"2591",-0.00183868646848162,-0.00337666806215886,-0.000588404066118819,-0.00614573865375911,-0.00545309353260282,-0.00260734410028152,-0.00160578748246154,-0.00831139764018973,-0.00887475166910923,-0.0174644522676406
"2592",0.00813916742933918,0.00774453861935531,0.00608333944796802,0.0123678736973216,-0.00387025132076557,-0.00224118023757935,0.000618675466692808,0.00392857545314884,0.00188939451517145,-0.00394991328905014
"2593",-0.00318682355154021,0.000240206699337886,0.00370573192434565,0,0,0.000467981741905321,-0.00395538773054238,-0.00495713260625308,0.00286978519899783,-0.00991407848530956
"2594",0.0109979171265011,0.0362543802514019,0.00699574292598681,0.0142529535675084,-0.00493797316119116,-0.002057812813263,-0.00868714629771594,0.00498182818920867,-0.00678599471483921,-0.00333780678179185
"2595",0.00581854585389441,0.008804599519183,0.00366648271958736,0.00878300148182709,-0.0120391347842984,-0.00515492010390906,0.00287918064186976,0.00417423993670774,-0.0101251479224939,0.00468855149106728
"2596",-0.000628745122446039,-0.00390450466222247,0.00115370877269672,-0.00373132486353323,0.00551664747226188,0.00263795526617727,-0.006615813408685,-0.003637485096051,0.00490641164241157,-0.00533332912498308
"2597",0.000838854255449606,0.000691722106677561,0.000768286737455437,-0.00124846019427671,-0.000327373381212359,0.000657297033333171,0.00113096163360926,0.00130403586810846,-0.00372390776974207,-0.00536192604130525
"2598",-0.00217933551447735,-0.00115225154362797,-0.00479765362783602,0.00149986317449247,0.00221145621925256,0.0010331152535128,-0.00928823272056845,-0.00572902641674378,0.00315639175310567,-0.0026954503170562
"2599",0.00252016083994944,0.00392161872353225,0.00385651947351207,0.00574129575770232,-0.00831315268470489,-0.00216080631199922,0.00608143426007679,0,-0.00910821418667418,0.00202706893995463
"2600",0.000377178644706211,0.00689343122385644,0.00307343225470258,0.00719812460873359,0.00512051902607724,0.00207164043791042,-0.00251899696725277,0.0112623911087262,-0.000167092841432237,-0.0107889326307644
"2601",-0.00121466236504353,-0.00251029368478695,0.00248938941791388,-0.00665363407292985,0.000657607928212123,-0.00206735761627297,-0.011993379696918,-0.00466206938085512,-0.0139573670880507,-0.00408999375384422
"2602",0.00117414188771248,0.0148709114647165,0.00248328866140568,-0.0111634550426732,-0.00492694626460954,-0.00225941090520265,-0.00434431234736921,-0.00208198761826828,-0.0100864720269586,-0.0239561487734999
"2603",0.00393716551600742,0.0114967139733668,0.00552595252273069,0.00827903301128208,0.000907825544999241,0.00018888002658346,0.00962541456891963,0.00573678089575491,0.00188373146773069,0.0140251252850372
"2604",-0.000167064293957742,-0.0104747010899641,0.000378997502040068,-0.0002488759122522,-0.00544159420872592,-0.00245301455182223,-0.00572020381311444,0,-0.00222204935950687,-0.00414932118355293
"2605",-0.000917892012507138,-0.000225274936745623,-0.00322029841756977,0.0126929322153517,-0.0000828203871567901,-0.00113510598651445,-0.00536961881358755,-0.00103690205051354,-0.00599569164882219,-0.00486111622344032
"2606",0.00179570830510123,0.00270318624579469,-0.00456093457862683,0.00663543504037478,-0.00116058466380475,-0.000378977041104567,0.0053986072767882,0.00103797833237484,-0.0000861869861390474,0.0160502406843015
"2607",-0.00204267667584068,-0.00292059213765783,-0.00267281621013316,0.00219727597498709,0,0.000758089907202164,-0.00536961881358755,0.000518451025256716,0.00396414164112247,0.0041208935885988
"2608",-0.00167091157220312,0.00788635845190555,0.00248843637359064,0.00414133392711813,0.00755287060539156,0.00511089625023642,-0.0026991377267167,0.00181417070636058,0.00283263519313293,0
"2609",0.00552350095021059,0.00581285024164857,0.0028643943677864,0.010189084106492,-0.002718489462054,-0.000658947345374861,0.00360881219901366,0.00517319030481045,0.00265340233410249,0.00547195189069516
"2610",-0.000915651883964252,0.0102243674701896,0.000761562717825015,0.000960889930470277,0.00371735676208074,0.00131923602314399,-0.00565042567954643,0.000257664187834683,0.00435379037351713,0.00136059565705837
"2611",-0.0177439957770149,-0.013861309470798,-0.001522167841016,-0.0170345972827883,0.014566539167425,0.00799911968082334,0.00529522923746795,-0.00360220305983294,0.0181895364523665,0.00679338516144568
"2612",0.00402844536462021,0.00133871228519755,0.00266772348384037,-0.0165978115266757,0.00113554297358398,-0.000280155263586379,0.00269774981410142,-0.00335632229531135,-0.00818100836312718,-0.00269901859172683
"2613",0.00650415311609387,0.0131462119588304,0.00817179520246158,0.0213453660160503,0.00234972075722673,-0.000280084378282308,0.00589357544765967,0.00595833480096908,0.00496594571106734,0.0196211203497609
"2614",0.00507734574318941,0.00241910355238284,-0.000565475745496147,0.000972017323326968,-0.00274819675406357,-0.00112102996159447,0.00292952236275923,0.00103055052736845,0.00418760461997314,0.00663567772410345
"2615",0.00221298537008119,-0.00153571227638605,0.00132023654526048,0.000971282898071024,-0.00672784001046278,-0.0026188051682221,0.00228605343757171,-0.00205841951537411,-0.00633864042804599,-0.00329593395865624
"2616",0.00233265775544167,0.00153807431599517,-0.00150689225782186,0.00388068155911903,0.00563080729545296,0.00206325388627548,0.00671566875312424,0.00386673419670092,0.00394495554763252,-0.00198416790706935
"2617",0.00477953586644109,-0.000877529086066087,0.0026409712969917,0.00483198284685571,0.000324554959557188,0.000561269388499985,0.00213983304453702,0.000256917626584974,-0.0010868489165885,-0.0218687617841493
"2618",-0.000206732632681228,-0.00483094027012687,0.000564411848504642,0.00360669644343625,0.00170354914339521,0.000654616516548634,-0.00615445077684862,0.00154036514386147,0.00887176074141882,0.00745254240077342
"2619",-0.00086880775946574,-0.00154454697821038,0.00206859494448941,-0.00527070787689443,0.00494015580207341,0.00252348130742841,-0.00391756333756244,0,-0.00331841709541714,-0.00806996786866232
"2620",-0.000248423243231377,0.00309384816061065,0,-0.00770704941389277,0.00249818651924483,0.000465880997370327,0.000253692749670575,0.00307648782469361,0.003995372099179,-0.0108473798076169
"2621",0.00795204159001139,0.00638909481232197,0.00900722161911238,0.00849499822094302,0.000104958596721438,-0.000522296990595916,0.00405895141346768,0.0091998899241359,0.000829033307186977,-0.00685405688185781
"2622",0.00332859823014475,0.00656747173922145,0.0210154936873836,0.00505428789671769,0.0118404232292375,0.00438823918094866,0.00985347772295841,0.00734359685123498,0.00737243201315074,-0.0048309230214546
"2623",-0.000737063303291485,-0.00587206797460693,-0.00382523307841043,-0.00119744113719622,-0.00620940360026556,-0.00167331412663807,-0.00312746676413667,-0.00276511091416909,0.000986777395059812,-0.00554777457712019
"2624",-0.00319699057409273,-0.00371914540978102,0.000731480962083308,0.000479586889692074,0.00544706251999361,0.00316606057000368,-0.00501954700284468,-0.0015124381856203,0.0112543741578648,0.00697340510093514
"2625",0.0018503008469033,-0.000219708449896827,-0.000365444120929537,-0.00119809526733772,-0.00478012086503288,-0.00185641829693661,0.00416227217488019,0.00403925731194343,-0.00528026816052429,-0.0138503695092584
"2626",0.0004923806066639,-0.00373365522887747,-0.00237616807229979,0.00599786911951328,-0.0026417553700282,-0.00158099878161133,-0.00163299069479927,-0.00402300735008854,-0.0065332382164125,0
"2627",-0.00151770118955719,-0.00286615495707809,-0.0089777447992917,-0.00763166332989051,-0.0015249374428904,-0.000931522115050987,0.00641607183180892,-0.00732143992050971,-0.00912454567818255,0.00561797306157019
"2628",-0.000205599148083158,-0.00508499718594435,0.00314299987707023,-0.00528717474433937,-0.000321680756951825,-0.000186482102597751,0.00662489456189097,0.000254311695897513,-0.00149328022653661,-0.0090782320655145
"2629",0.0048900788276911,0.00577767753859493,0.00552887086389786,0.00483198284685571,0.000160922477482117,0.000373182712740672,0.00211103795666023,0.00991606467621819,0.000997025581613187,0.00422841721504996
"2630",-0.00126766300448045,-0.001767589169265,-0.000549748065779343,-0.000240394564499979,0.0154365460168222,0.00521979004746975,0.00322174503483996,0.00251790216787939,-0.00547811241339369,-0.0175439077995795
"2631",-0.00192438099687786,-0.0099601816346705,-0.00971938998542299,-0.010341604739158,-0.00158336268466253,-0.00176178525729531,0.00345870454507846,-0.00502300476757667,-0.00417292605575026,0.00428580271427803
"2632",0.000218609436818173,0.011178202693789,0.00407407114701863,0.00170120067964152,0.00198220960001372,0.000557409592365277,-0.000615484160056301,0.00349131064587405,0.000167582970164393,0.00426729339038379
"2633",0.00832502448285166,0.00375881087762608,0.00313530734976752,0.00994653172067128,-0.00142446786413108,-0.00278525803045782,0.00172417644953904,-0.00126985101630639,-0.00762523906905432,-0.00637392368741607
"2634",-0.00674415191930677,-0.0104542114958639,0.000333111038648415,-0.0110526289881859,0.00895626033597807,0.00251363547711336,-0.00331986543389717,-0.0162723550814567,-0.00211095161698893,-0.00997862781066583
"2635",-0.000246885416969711,0.000226749285485051,-0.00147982532957791,0.00219626531679329,0.0020422882968798,-0.0000927191450764697,-0.00394747006812257,-0.00258496419557419,0.00287694195295307,-0.010799137029343
"2636",-0.000452740876513147,-0.000906545544664628,0.00203784116627848,0.00511309246370284,0.00219527340440506,0.000928760912779936,0.0019815571716848,-0.00414584276525587,0.00337496633584977,0.00145565913800816
"2637",0.00119439226514451,0.00340291356901368,-0.000739550872532968,0.00532946491185071,-0.000469305182578816,0.000278241285447844,0.00395527673638663,0.004423537632122,0.00428861426654237,0.00436033063266361
"2638",0.000657977673661048,0.00339129940839777,-0.00277520282814159,0.00963865245639139,0.00375612832998162,0.000834946053343888,0.0064025557874472,-0.00207260097979423,-0.00895921460269622,0.00217088652750053
"2639",-0.00805611153481089,0.00247857837845089,-0.00241184708659115,-0.0116945749904104,-0.0106813004829386,-0.00491242536787651,-0.00591217962831658,-0.00519231055488978,0.00380193474314017,0.0115524115461247
"2640",0.00895029166053996,0.00741739943785169,0.00446332153285911,0.00772768572641791,-0.00330977446775116,-0.000931522115050987,0.00136561621971154,0.00104401347255623,0.000757545673891968,0.00642396808240298
"2641",-0.0087888956557215,-0.0111556618587599,-0.00999808360810484,-0.0127005476569155,-0.00838173574823986,-0.00372910595561837,-0.010911258554913,-0.00469220913040413,-0.00487806551929248,0.00425518775965816
"2642",0.00186445972132443,0,0.00336643031363892,0.00461158943426732,-0.00231213758538684,-0.00233962192027848,0,-0.00209536914389596,-0.00253552231237308,0.0204803110442378
"2643",0.00169570953440989,0.000451178307552702,-0.00484619131599373,0.00579841472163212,-0.00321966590027156,-0.00367304491615028,0.0106558058722537,-0.00892408081069085,-0.0163531693701027,0.0103806233302839
"2644",0.00231202953846799,0,0.000187203399183433,-0.00192173108050331,0.000240994967753982,0.000754526202326744,-0.0112874925618164,-0.00158875351704613,0.00370403148260934,-0.015068498558463
"2645",-0.00914440322625842,-0.00360853298729791,-0.0073033886418894,-0.0120336868819894,-0.00827388975647569,-0.00188447256931767,-0.0174381848549621,-0.00503986300930548,-0.000429076564428699,0.000695472358283933
"2646",0.00648505774827424,0.00203709259007967,-0.000565914028069936,0.00194888349531563,-0.00599371858466624,-0.00160479281419912,0.00485161228517517,-0.00106658976957175,-0.0102172404033893,-0.00972898790088284
"2647",0.0010739556867907,0.00225900363642517,-0.00264238117730253,0.00948214437756212,0.00146693640063011,0.00132344813986851,-0.0073697134987335,0.00186815765733783,0.00164817836266629,0.00421046853524154
"2648",-0.000742752349902398,0.00135220535832192,0.00681289532439622,0.00818873633241224,0.00170863149065936,0.00132208043181503,-0.0011520332402617,-0.0061266042863749,0.00129905602061964,0.00978337842656662
"2649",0.00751481141276544,0.00855292376686734,0.00695488342600692,0.0193502599112181,0.00690428466771476,0.00292323263158778,0.0125594606462391,0.00696861741539623,0.00354606460267948,-0.00484429563586741
"2650",0.00168022055275197,0.00423996572647556,-0.00130662967050288,0.00492156787414322,-0.0062922889559418,-0.00103436721303651,0.000379647791835858,0.00452505051216945,-0.00180986815314899,-0.000695400785539535
"2651",0.00466406691502375,0.00622222942524431,0.00242987953736984,0.0125932445211472,0.00121761836227607,0.00141191665421703,0.0101212720009614,0.0135132387643344,0.00820235710585404,0.0111342268915033
"2652",-0.000122230135127133,-0.00154589623009171,-0.00130524626281836,-0.00460611970031621,0.00275695012929544,0.00122159739831185,0.00400816626741629,-0.00235275774854049,0.00445323296531375,-0.00344110942841314
"2653",0.000529565466281356,-0.000884784996381782,0.00522774969351603,0.0030077800777697,0.00873303172459639,0.00366133880157893,-0.00249491576460226,0.00943385247189577,0.00699121828807892,0.00414366093869045
"2654",0.00541390186871915,0.00199237302958721,0.00408620228002854,0.00830454740557163,0.000400859631271233,0,0.00800375743846371,0.00700935821029058,-0.000253992039166984,0.00894087224434292
"2655",0.000445400031027221,0.00552378588307523,0.00369965090945601,-0.00114387764377555,0.00288456041696428,0.000280343228975743,-0.00397016509183445,0.00438263882764089,0.00135497965184661,-0.00136337802319941
"2656",-0.000890136550733667,-0.00593265522974351,0.00184298758060231,-0.000687191244042262,0.00423459622512778,0.00177652063361178,0.00211754469803971,-0.000256800260155288,0.00862655630288489,-0.0136518315761254
"2657",-0.000243148854322195,-0.00309474152784972,-0.002023595660401,0.00297963861122863,-0.00389848661980186,-0.000653485853657321,-0.00261031278145962,0.000256866223468322,0.000419218507140329,0.00207609617564697
"2658",0.00243082996150035,0.00221723722183498,-0.00350232201257372,-0.00251361618766954,-0.0130193319266865,-0.00560378835679831,0.00124632523659129,-0.00154009488397822,-0.00326879562934856,0.0110497861959944
"2659",0.0000405460129913049,0.00774344997633891,0.00332961185741221,0.00824727354006116,0.00161859367076045,0.00319353917765053,0.00535231981102369,0.00437021493744671,0.00807264561171617,0.00956278073642225
"2660",-0.000929695711457401,-0.00461034122648374,0.0033186399283438,-0.00545324891574994,-0.00492850793558508,-0.00159149235970879,0.000866551305555019,0.00179171353858809,-0.000750717402837386,0.0060892964033703
"2661",-0.00117293022230147,0.00110275031001827,0.00294005249948737,-0.0004570415748405,0.00592719573402722,0.00168774229956914,-0.00210297227577405,0.00383242325680166,0.00751315629423854,0.005379955507687
"2662",-0.000567106055553657,0.00264380496933381,0.003297889678332,0.00114293008532473,0.00121084008916839,0.000280755056114357,-0.00012373374263841,0.00152682426159512,0.000497124857119502,0.00602005367344782
"2663",0.00222878698736273,0.00483419113356365,0.00584376925547625,0.00296797574029717,0.00702100955407436,0.00248424258468782,0.00446304854885615,0.00330379597043007,-0.000828140786749532,-0.011303174426881
"2664",0.000485234741016249,0.00109315572547009,-0.000544798787692202,0.000910509621702582,0.000561474667140072,-0.000935135190454073,-0.0062946942142591,-0.00253278438853488,-0.0020721093730276,0.00201745736003356
"2665",-0.00193980413974471,0.00152913090020013,0.00254317493248379,-0.00409361489783533,0.0103440050502126,0.00346288509474735,-0.00347771690112297,0.00126948624761236,0.00157802322960099,-0.0073824498756202
"2666",0.00182203709220263,0.00196298990836996,-0.00090596590559755,0.00365397635315112,-0.00849211598888622,-0.00270497199723163,0.00336521946130564,-0.00202897309091632,-0.00779495838112476,0.00202830017005384
"2667",0.00185921076206674,0.00108834778293976,-0.000362657722954074,0.0068257863365071,0.00112060064648389,0.000561049209975684,0.00074535216977889,-0.00355795986248686,-0.00117007937868652,0.00202433339157682
"2668",-0.00246087657747307,-0.00652317620356047,-0.0010885014979255,0.000225896354356436,-0.00359791355675143,-0.000840829044598257,-0.00546182650051696,-0.00382533868860191,0.00292861680313594,0.000673322171594659
"2669",-0.0000405034063132304,-0.00131311597442085,-0.00617517044834115,-0.00903733055323575,0.00545674844884569,0.0012159821510298,-0.00174737136132797,0,0.0120974218913947,0.00672959153000807
"2670",-0.0141152128583242,-0.0149025633007289,-0.0104165090314569,-0.0237118607327462,0.0085394195945363,0.00373713023728772,-0.00762681103099605,-0.00972852474530506,0.00741901751576979,-0.015374396255745
"2671",0.00147676769327254,-0.00200222091806601,-0.00147752107875521,0.00233523028956384,0.000474907355218379,0.0011171031752224,-0.00478763987141884,0,0.00474594554247565,0.00339445675241579
"2672",0.0099131155002905,0.00735612480624503,0.00739781687360686,0.0102518200426747,-0.00514132467429351,-0.00241765156599572,0.0153183187589956,0.0067216116864699,-0.00708529190418361,-0.00879568904694039
"2673",-0.00012147674399976,-0.0011064108064659,-0.00128505974759974,0.0011531108813676,-0.00421356468750445,-0.00298229155115493,-0.00286800500426643,-0.00487891477338764,-0.00770993286925747,-0.00477816212774163
"2674",0.00174417036498942,0.0053169668268096,0.00330880174144288,0.0103662920402989,0.00367266239570685,0.00186969247874358,0.00437683827263102,0.00851585398150445,0.00735658768333813,-0.00274344684758798
"2675",-0.0155907485836809,-0.0125605822554546,-0.00677911325998404,-0.0127679909094521,0.00747748052191111,0.00354565046895594,-0.00684780766035453,-0.00639713899049277,0.0050873470479853,0.00275099405355195
"2676",-0.00156310747418342,0.000669354823279678,0.00442732811660407,0.0085448900780305,-0.000237093989575943,0.000186086333161084,-0.00739621192947681,0.0038631434876979,-0.0015511062380783,0.0178326868731391
"2677",0.000782711555319393,0.000892182691481613,-0.00220379069623278,0.00366394377781876,0.00244842972684167,0.000650470417126625,0.0089670900675074,-0.000256545660889618,0.0037612345765845,-0.0121294223954782
"2678",0.0104569738532776,0.00579305090218196,0.0020246161845503,0.0111796189531808,-0.0038602938440051,-0.00195090216563976,-0.00087619389582283,0.00179618830258299,-0.00448031110328595,0.00272854600406491
"2679",-0.00358543352193563,-0.000221407049130096,0.000367398123751084,0.00473824451008187,0.00680154929985277,0.00344417993692581,0.00826842787056647,-0.00076857684043663,0.00376400461307602,0.00884355670473025
"2680",-0.00233063331398342,-0.00132950601562642,-0.00514151080280079,0.0031439892039391,-0.00369207682876316,-0.00157699221605001,-0.000994017674374348,-0.00358847897656034,-0.00309771750383503,-0.00067436901525264
"2681",0.00233607785485601,0.00710000197454397,0.0033223928849313,0.00582034168804002,0.00386339678776171,0.00167226965114353,0.00472641687584097,-0.00128638896933564,0.00367975301594758,-0.00202419449601332
"2682",0.0000410201763978435,0.000220450578507059,0.00110371962339451,-0.00356097825208868,-0.000628268700106793,0.000927754651473656,-0.0050755121707966,0.00309083528100529,0.0158872741712119,0.000676053664256049
"2683",0.00114472916204078,-0.00396482145179744,-0.00202144197934651,-0.00178704390292839,0.00322229259311113,0.00231665636089518,-0.00149312942444191,-0.00205428961222842,-0.0021654021627171,0
"2684",0.00473761952962448,-0.00176925059317024,-0.000552367964517964,0.00156635465210631,-0.000313385296431545,-0.000832116178486886,0.00535833613856695,-0.00154393501013506,-0.000482213478254612,-0.00743240066882345
"2685",0.00601615452527926,0.00731076026477973,0.00792194705362803,0.00156402494620855,0.00297783280523545,0.0015729835753544,0.00644504924390099,0.0108247815007008,0.0117401012243479,0.0279101820157066
"2686",0.00141417394267718,0.00219909935644313,-0.00402114642522244,0.00736112729552696,-0.00764902160033309,-0.00294234604378707,0.000123035725395848,-0.00382460609005097,0.00190747099030353,0.00132448516535044
"2687",-0.00718211453977613,-0.00636381355168492,-0.00440450025395356,-0.0130647164839849,0.0158578384350643,0.00696011788022766,-0.00209308984444356,-0.0010236043299422,0.0111058307330769,0.00198403176737982
"2688",0.00341371645766619,0.00706709800346461,0.00423953659091159,0.00650673028216286,-0.00613532257135019,-0.00239632935809686,0.00197420143595162,0.00614899246527667,-0.00509964698807197,0.00990112731437764
"2689",-0.000121433187195819,0.00899132801944358,0.00587372632715555,0.00735603676465235,0.0102367133158339,0.00434200897551817,0.0065272233463276,0.00814865284864807,0.01040932908145,-0.000653653071059468
"2690",-0.00117476519013726,0.000217385571476214,0.00310226346515519,-0.00663858559987907,-0.00216569787328769,-0.00073591542621787,-0.000611692910802208,0.000505215887647514,-0.00124876292637321,-0.0111183607233376
"2691",0.0106658834718754,0.00760530850746077,0.00454793933934505,0.013366093206266,-0.0119380876132479,-0.00570709111154133,0.00844748773863158,-0.000252707043361333,-0.0139095021183909,0.00198403176737982
"2692",0.00337088775935879,0.00452874261970249,0.000724245543419322,-0.00109914189571647,-0.00525661094640351,-0.00240688623292173,-0.0100763659797605,-0.00429287365259745,0.00293205479147218,0.00264029608816352
"2693",0.000479677448728566,-0.00601119396151795,-0.00199048611689334,-0.00528163444534879,-0.00394338779781334,-0.00204128044881879,-0.00367924126320218,-0.0073546138152264,-0.00750629752696419,0.00460829992672163
"2694",-0.000319696849482409,0.00323984435208113,0.000181305514558971,0.00265470848013249,0.0041173766223892,0.000185825073726553,0.00615435739497383,0.00204391421407935,0.00437865612309007,0.000655366512221311
"2695",0.00134605299396728,0.000430582663460077,0.00145044824493246,0.00595771155445157,0.000394289254649349,0.00120859452573652,0.00415964899971488,0.00324024336909634,-0.0049936983197939,0.00458415661069123
"2696",0.00212701246829172,0.00193672965234049,0.000180857721601813,0.00350961454005239,-0.0057544099768353,-0.00390024834303448,-0.00536069570078979,-0.00281964803228241,-0.00932046530168462,-0.00130376311982083
"2697",0.00100102908307731,0.00472507943253531,0.00579192340438883,0.00218567337949183,-0.00245787654382401,-0.00111851808276509,-0.00771657539844384,-0.00308481050558718,0.00209072047209125,-0.00195826488688433
"2698",0.000360115112502113,-0.00299270043527522,0.000359927205674015,-0.00458013104452448,0.000715592917668761,-0.00195983839467706,-0.00246905350490745,-0.00257884422901922,-0.00802439396506838,0.00850230752397341
"2699",-0.00267932367874169,0.000857564043424519,-0.00395754761854195,0,-0.000556158202328239,-0.00130900565419512,-0.0032173411737576,-0.00698014871686758,-0.00760397166468274,-0.00389106408858941
"2700",0.000200457998094095,0.00214228238724612,0.00108366283358574,-0.00569671116505566,0.00286074162232453,0.00177891983665934,-0.0059589231497913,0.00442577488138074,0.0045647049233779,0.0039062636106455
"2701",-0.00204458347217285,-0.00769565128829386,0.0021649036297271,-0.0169678957891104,0.00625997465094885,0.00299079431004712,0.00537027034841708,-0.00544304218010849,0.0104673890046638,0.0168611887231829
"2702",0.000602612874618158,-0.00301590982561017,0,-0.00268981929711609,-0.00181114794649639,-0.000838430094397991,0.000275519929850754,-0.00208497785656325,-0.0111619690930858,-0.00892858080554015
"2703",0.00389436948612487,0.00172856351545803,0.00198001862051678,-0.00359638814911922,-0.0150679613252256,-0.00512999868539643,-0.00801607644832159,-0.00443989301806158,-0.00942013975491429,-0.00386108364400783
"2704",0.00119963682591218,0.0034512082986311,0.000718747222891114,-0.000676901962286758,-0.00296330054367988,-0.000187410293433166,0.00744964730175179,-0.000262358724170242,0.00188552217038396,0
"2705",0.00351524008555537,0.00752382400794294,0.000179496355366515,0.0115125349491563,0.00224900982528453,-0.0012191357256236,0.00112786311863555,0.00708467255114398,-0.005155036454914,-0.00516788856168493
"2706",0.00433855230449254,-0.00192027048789634,0,0.00022316911304987,-0.00183100940521685,-0.0011374894948859,-0.00200284641327342,-0.00234476912830739,-0.00666232099584918,-0.00844151018349193
"2707",0.00214005912307647,0.00320650783702958,0.00592365766884351,0.0158409447401351,0.000965727696105478,0.00141203383672672,0.000752495132553932,0.00470080794361638,0.000496853535568054,0.000654869887072751
"2708",0.00118656096045888,-0.0017046915126967,0.000178350991032694,-0.000219474960154287,0.0000801303566109191,-0.000281897135988807,0.00639260206200798,-0.00519888074226238,0.00281383757653186,0.00130894998339981
"2709",0.00592507102839201,-0.00128062655006633,-0.0005352203767226,0.00746925832899636,-0.00377774519039598,-0.00103439196291288,0.00311367813824548,-0.00130659011641931,-0.0053643724579413,0.0111110931727056
"2710",-0.00113872162183504,-0.000854977207798147,-0.000535506990976042,-0.00501527458137319,-0.00282389213979284,-0.00122341298252271,-0.00360068329900742,-0.00183114735350287,0.00472949729661876,-0.0155139513659167
"2711",-0.00165113331219713,-0.000427819587952682,0.00125022964475496,-0.000657428830499796,0.00315563588830248,0.00113062697797628,0.00199383200063652,0.000261903496820759,0.00817578687507758,0.000656522276818006
"2712",0.00263828581651726,0.0106997654798837,0.00713519239195093,0.00986843785797809,0.00161319347999656,0.00037663268560606,0.001367855249365,0.00707548306739159,0.00262123193608743,0.0118111334310549
"2713",0.00157097348150548,0.00254071499864006,0.00513633151705339,0.00456023874660083,0.00193253696498186,0.00112915397177615,0.00422253201278511,0.00572452952935776,0.00318626628780616,0.00194549867153038
"2714",-0.00149009803831268,-0.00190064406309676,-0.00123341239342878,-0.000432371150681843,0.00425978760228451,0.000939897035002524,0.00655471589460066,0.000517614316628112,0.00081438227205477,-0.00129448070386373
"2715",0.00121740592952713,0.00169281124954779,0.0123499498230846,0.00908309484126502,0.00720280211503965,0.00338024532941605,0.00221138217905326,0.00284468469636345,0.00756775170939661,0.00972125587305173
"2716",0.00133370369932084,-0.00253490279838853,0.00453129240213035,-0.000642916334573029,-0.000715081699876774,-0.00168434964210684,-0.00502607471162453,-0.00128931500312801,-0.00686479567113552,0.0025674912770961
"2717",0.000704968219083391,-0.00381200579917451,-0.00104098559974786,-0.0051470079022089,0.00127239561106451,-0.000375079158876912,0.000862447681811984,-0.00103275294311445,-0.00683096684694662,-0.00128045807361343
"2718",0.000978560524540262,0.00425177489707229,-0.00104192419119808,0.00237120384757872,-0.00659167986447839,-0.00253194026611225,-0.00110818127414281,0.00439374532233971,-0.00376647024727261,-0.000641082861988718
"2719",0.000273820985131623,-0.00169352791643484,-0.00226007652588278,-0.00881715724765808,0.00175883688991396,0.00103437443437082,-0.000739339765497338,-0.0012867524841671,0.00591765440811454,-0.00448993064839287
"2720",0.00516049770534766,-0.00296865540720381,0.00226519604228437,0.00368844251210443,-0.0106136061898209,-0.00413236757083402,-0.00320686089460276,-0.0043801609575671,-0.00637305340610395,0.0051545684159735
"2721",-0.00388946797575207,-0.00318997985290459,0.00243389338814159,-0.00799832092118014,0.00177452317683024,0.000942848342256664,-0.00470169856922187,-0.00879923091807633,0.00156238794866881,0
"2722",0.00175703213368217,-0.000640213656170174,0.0083246310487417,0,-0.00619968733357668,-0.00301488298937269,-0.00497269670440581,0.00156659935921799,-0.00385879300840419,0.0102564681117521
"2723",-0.00494996046314744,-0.00106734332578851,-0.00808394038986626,-0.00217902904913525,-0.00478030724294742,-0.00160635183832347,-0.00387322132119738,-0.00782062106895687,0.000164806722742883,0.00126895282363715
"2724",0.00129250600658537,-0.0023510075630726,0.00537531157127957,-0.00677008381689237,-0.00333759963052993,-0.00132522504801669,-0.00614548454379149,-0.00157644681933555,-0.00840540598937634,0.00443606490635928
"2725",0.00817612056139683,-0.0017138445092274,0.00758882696244489,0.0145117738545222,0.00661620313773481,0.0032225440448177,0.00454319788314583,0.00447362056416933,0.00473697324462785,0.00504724945748625
"2726",-0.00372497273609707,0.00579414385563082,-0.000342224216783982,-0.00628516408385671,0.00957468630022484,0.00358990293015826,0.0021354039360082,0.00104815353069121,0.00190235728862942,0.00251101593966951
"2727",0.00155781695008894,0.00512055149744217,0.00428082565078625,0.0093782988984481,0.00032158712207786,-0.000658840371598579,0.00188048796883034,0.00680426478035256,-0.00379756469406989,0.00250479097826695
"2728",0.00132222768613621,-0.000849169652790027,0.00562657321151661,0.00518595723478743,0.00445229461229446,0.000603510957974729,0.00075083303778567,-0.00441899618615471,0.00364633303466189,0.000624536740310377
"2729",0.000388493293851377,0.00254935127104194,0.0011867955336029,0.00128986392146779,0.00440913373512797,0.00132034488674293,0.00625149361227351,0.00391626599708772,0.000660564770369465,0.0062422403245177
"2730",0.00333861555962334,-0.00254286860572972,0.00237088435130262,-0.00515246354835497,0.00271334242234222,0.00160063870310556,-0.000621153130118679,0.00130038100577012,-0.00470335003377598,0.00620332494232834
"2731",0.00154750865454401,0.00212453240527521,-0.000168841665999064,0.0112213387505851,0.00374101762670143,0.00122227097657346,0.0115628674393815,0.000260108352175381,0.00853920555780463,0.0191123283471131
"2732",-0.000695211506337334,-0.00826798166832587,0.00794185887591392,-0.0064019070598369,0.00420253507130308,0.000375360919094625,0.00712878605920375,-0.00259680144991647,-0.00361695842799903,-0.00604964843524292
"2733",0.00170080643271864,0.000641167009796328,0.00620272249560827,0.0047249069472235,-0.00221090892106024,-0.00122002321212356,0.00671225878703452,0.0093723981910796,0.00346504416685955,-0.00182590324516907
"2734",-0.00362761148428892,-0.00704959311855169,-0.00833047684811195,-0.006199061422417,-0.00284892598955488,-0.000375976357178121,-0.000363613270441543,-0.00232142717752781,0.00411082802213669,0.00182924326638534
"2735",-0.000310072765576597,-0.00150607821477788,-0.00739249307729961,-0.00430213562601367,-0.0150795263379195,-0.00507690931281679,0.000606238096099165,-0.00180949318266743,-0.00818799659841141,-0.00182590324516907
"2736",0.000930076156683723,-0.00452483926223912,-0.00440076371327214,-0.00216029240713156,0.00209518971187195,-0.000472284154907077,0.00363598681603339,-0.0049211226106739,0.00148601506198331,-0.00304873877730882
"2737",-0.00232256060368319,0.00216435176212992,-0.00527036078783605,-0.00671136322344401,0.00675451837457475,0.00141819131074294,-0.00157007935423981,0.000780652350691247,0.0020608359090073,-0.0134557875869372
"2738",-0.00500526884239572,-0.00453549612363968,-0.00734920861565369,-0.00523107598471484,0.0108627637774783,0.00358713723395065,-0.00858721672371965,-0.00130013407844909,-0.00123390920095268,-0.00123984494504614
"2739",0.00850087718323467,0.0065090463780475,0.0154959112626565,0.0208150844069814,-0.00869162692892445,-0.00253959433452089,0.00670991029651291,0.00937474647342129,-0.0000823820086522931,-0.00310368377575998
"2740",-0.00293871198830109,-0.00129341861017118,-0.00491699959678382,0.00493660007002217,0.00741236956370872,0.0013201351181642,-0.00460483762538466,-0.000257781793636336,0.0120263507079679,0.0161893255167598
"2741",0.00170639982593501,0,0.00494129594696258,0.00512614452943461,-0.000395376058591856,-0.00160109975107436,-0.00206988132840635,0.00258047337375955,-0.0126160099901025,-0.0079657033931777
"2742",0.00654275482771904,0.00539595439870277,0.0091556570158946,0.0133870097920681,0.00316611745258033,0.000188852056335564,0.0071977946453945,0.00592028633606212,0.0016487017005804,0.0067942881877463
"2743",-0.000884513486821281,0.00364965680509344,0.000672011076320755,0.00251643847575145,0.00323506410967922,0.00320656969433619,-0.00278585493357508,0.00230276962497822,0.00921730706580015,0.00552146022906941
"2744",0.00230958724768371,0.00919797024688762,0.00822700480133265,-0.00209167843817271,-0.00275260751857831,-0.000846153208006739,0.00206499772646707,0.00459547319545628,-0.00252790514216528,0.00305072465542766
"2745",-0.000499041597079475,-0.00635873670484333,-0.00432969481574852,-0.0146720340597649,-0.00141971349141057,0.000658656615743825,-0.00412149796755046,-0.00101648109042951,0.00416940810987576,-0.0018248551037251
"2746",0.0101447701992508,0.00639942898884471,0.00301051699395227,0.00744533397982883,0.0013427178112777,0.000188089287598725,-0.00219055032780457,0.00432468941900233,-0.000162859233691082,-0.004265696046719
"2747",-0.000608816041584248,-0.00402725512001911,-0.00200101071674508,-0.015836182425789,-0.00985910467615758,-0.00319632046998375,-0.0012200059062667,-0.00658553559365116,-0.00626982340639715,-0.00673198010526599
"2748",0.00875513193564603,0.0010640516553877,0.00100247623338268,-0.010941947097166,-0.00334535866585428,-0.00311259007986908,0.001099182164227,0.00484437140640726,-0.00770241717713527,-0.00431300522668032
"2749",-0.00207543388104936,-0.00361380563453839,-0.00450676576878439,-0.00563989118715535,0.013494578315842,0.00369555546521627,0.00183001713099307,0,0.00404622632611429,0.00866337563776698
"2750",-0.00121013120178581,-0.00149363890574383,-0.0105633464877575,0.00196348538738667,0.000473994488235485,-0.000471811240758346,-0.00767176065739106,-0.00380608318027376,-0.00337195504143284,-0.0122698975885782
"2751",-0.00359650332582628,-0.00363240756206962,0.00254186589807004,-0.000653204764547444,0.00497604331310852,0.000755340031078244,-0.00589027515281237,0.00382062479604817,-0.00709688067337855,0
"2752",0.000189947272477564,-0.00171568216729523,-0.00371865925582493,-0.0135076482232015,0.00345813654853577,0.00207609281032028,-0.000370256271098879,0.00177621631805036,-0.00207779255319152,-0.0167702126206949
"2753",0.00315301409855606,0.00257792287302783,0.00644721395235592,0.00287089468958812,-0.0078321788075032,-0.00178936534186547,0.00407528106125254,0.000759572353670634,-0.0131590072457732,0.00315851657128929
"2754",0.00545328655894894,0.00514240251525622,0.0047200619510237,0.0116714691581135,0.0000790090676017208,-0.000754695754718204,0.00332044485937821,0.00379678147675255,-0.000084353111390878,0.0050378444325565
"2755",0.00301283926526685,0.0019187490651893,0.00335584587284732,0.00500663473453589,-0.00205247660159025,-0.000660943464963593,0.00110302128772677,-0.00176490012569663,-0.00396692258692799,0.00250629588749507
"2756",0.0017648269973467,0.000425359164795136,0.00183942148337168,-0.00671436306478779,-0.000395540210436307,-0.000850468972762419,0.00404064858220377,0.00303095653149876,0.00118634012056029,-0.00875007309041997
"2757",-0.000112253789080197,0.00212679172231534,0.00400609987981526,0.0119931079624347,0.00751736154553417,0.00406618625384358,0.00207341591939869,0.0095696085028385,0.0086330595237738,-0.00441362391405054
"2758",-0.00408624663726131,-0.00594230491781478,-0.00465507011993149,-0.00732611290316565,0.00424099646642162,-0.000376677633114109,-0.000608592459913404,0.000249229701419162,-0.00201391293134034,0.003166583158283
"2759",0.00832738697297053,-0.00106734332578851,0.000501070664865377,0.00217067846384533,0.00375373519930444,-0.000188255690238504,0.00414036858022437,-0.000727081656357709,0.00210207685192976,0
"2760",0.00634127444789301,0.0132506506673211,0.0120200245679378,0.0112626562956981,-0.00911581046115273,-0.00226141275130542,0.00557837238702796,0.00978431572030947,0.00461489343849641,0.00441919659547785
"2761",-0.00384047830344925,-0.00105460237564581,-0.0101459996331033,-0.00528345872643632,-0.0129737073168493,-0.00453382411682479,-0.0192564283156933,-0.00322971950847373,0.000751666230226267,0.00754251726589228
"2762",-0.00052391085768555,-0.00401183437403563,0.0013420328098912,0.00131148004809045,-0.011073115848839,-0.00294099287768179,-0.0104387539157925,-0.00174504740838666,0.00267066432982821,0.0056144599261303
"2763",0.00205966748022623,0.00420363536635415,0.000670082062594002,0.00654881160469367,0.00582843738314653,0.000705541764169482,-0.00364200185720243,0.000749450115848482,0.00141500750303813,0.000620211184653829
"2764",-0.000261554027750743,0.000849946530373957,0.00468787097035905,0.00845801894307985,0.0013642969770975,0.000380546937438497,0.00630204486791452,-0.000499200331025018,0.00523650578067514,0.00433987205688369
"2765",-0.00119637588567412,0,0.000499868570691397,-0.000860263571421882,0.00296547550007165,0.000381014013626668,0.00488501495226212,0.00149784798730468,0.00686286577041728,0.0148148021084444
"2766",0.00048658289565795,0.00148621768484358,-0.00133242132905464,0.00258296726160245,0.0130253513578409,0.00428232115805471,0.00361423405380035,0.00648069247049876,0.00377766289999992,0.00243299406141095
"2767",0.00205749630382535,0.00233197659474516,-0.0023348396111762,0.00686985699802434,-0.000867622066221707,-0.0012321788640387,0.00583715812402286,0.00346692055979458,0.00507236345236772,0.00485430284159838
"2768",-0.00377051868079681,-0.000422961613844808,0.0018388476075053,0.00469091570300351,0.00157891561900358,0.0016131018532124,0.000246972031916703,-0.000740436398890876,0.0065120391780551,0.00301940706457482
"2769",0.00715725319849669,0.00677113914273342,0.0060069531888074,0.0188878983118048,-0.010799138058993,-0.00331526673851235,-0.0050609691767427,0.0059273264347337,0.0121310147653697,0.00481637198410567
"2770",0.00632496389842396,0.00273217623081679,0.0137668217093292,0.00958134854019654,0.00478123963795918,0.00104528261661163,-0.00161284861879629,0.00564692826249846,-0.00263685173572759,0.00599165342118746
"2771",0.0042148977141967,0.0121567598871897,0.0122709073735359,0.00495153357925626,-0.000158801660173014,-0.00047443865236263,-0.0156583953797973,-0.00146470578995284,0.0051273754206056,-0.00119116894609306
"2772",0.00666424689832734,0.00683369380954124,0.00274773656383176,0.00862248921879472,-0.00285541151590063,-0.00123479449748187,0.00101034986087245,0.00440093813557363,-0.00103616292871167,-0.00357789130999808
"2773",0.001828623554889,-0.00267366770619726,0.00580278972771398,0,-0.000636467516198835,-0.000475791747737597,0.00567531525579046,0.00024323687121508,-0.000159610625395157,-0.000598312713800175
"2774",0.00226342190109041,0.00144352502678902,0.000640913644922581,-0.00162838161748524,-0.0133724187532713,-0.00475728528383401,-0.0115376381694333,0.00146021556165055,-0.00462848144008432,0.00658673582176394
"2775",-0.00152989246782176,-0.00329494544409104,0.00640611950100123,-0.00632010348777057,-0.00121017367793308,-0.000286406074842538,-0.0121795611084948,-0.00680409737667242,0.00240516309456029,0.00356925525226215
"2776",0.00729594353335883,0.00702491688845797,0.00668363026731567,0.00615513024182257,0.00411954500993961,0.000669133900198071,-0.0034679938025397,-0.00122341539773729,0.00327923700935173,-0.000592638145727076
"2777",0.00651907720624578,0.0133358879511192,0.00316161496525735,0.00958393850193828,0.00168910075548068,-0.000668686459419421,-0.00811937711020372,0.00710420607012918,0.012117322829762,0.00652416725529137
"2778",-0.00341820123719605,-0.000809784388957513,0,-0.00383747265119616,0.00417638810799126,0.000477654847991227,0.00272869405089349,0.00316227042855455,0.0016540564087435,-0.00471419813690632
"2779",0.00953154129153244,0.00445792620218222,0.00803659223518749,0.0131791967949453,-0.00135975933893773,-0.0021983546081259,0.00712704433370237,0.00703219923095966,-0.00809938677517319,0.00118411653188644
"2780",-0.00168066831868086,0.00100865265717176,-0.00844144502725697,0.00120063992084551,-0.00928964392021281,-0.00316117470535016,-0.00977862021551723,-0.00120408638914771,-0.00221973998905778,0
"2781",0.00454950508340857,0.00483685850673776,0.00630613394398227,0.00819500618930746,-0.00525426848602095,-0.00259463519578584,0.00649703512955147,0.00120553796099809,0.00444936433776144,-0.00177407408737407
"2782",0.00813085776362521,0.00681912623287406,0.00422993907131608,0.00574948886583337,0.000975000989480668,-0.000385369292986271,0.00813311338174216,0.00650109431775991,0.0018193640534625,0.00236963602636964
"2783",0.00212282665788099,0.00298793951850596,0.00608427776164944,0.00473094511189354,0.0043028253973969,0.00289168859280031,0.0138301249324346,0.00406721925048203,0.00497431496290068,0.00709240651970733
"2784",-0.000388697909626701,0.00317763517712466,0.000310144382704935,0.00843638542871394,-0.00541598783661601,-0.00192210226126344,-0.00353661094438074,0.00619471941448357,0.0121778992157284,0.0105631140112774
"2785",0.000423920707893544,-0.00395948359142995,-0.00480551250995565,-0.000583783052441111,0.0082086785942066,0.00221458261850915,-0.00190146527998114,-0.00331515525623938,-0.00667547144802505,-0.00580700294982217
"2786",0.0115777342394479,0.00795061829784083,0.0073208844573267,0.0138214077451466,-0.00370817745763197,-0.00297851292678541,0.000380953780398929,0.00855310771589934,0.000781480028276382,0.00759347409706135
"2787",-0.00662981797029683,-0.00985990198654518,-0.00850464157701281,-0.0151690234855846,-0.00695857857447768,-0.0025055252934596,-0.0128219363775774,-0.0150764929320545,-0.00562199547627107,-0.0028985109481735
"2788",-0.010257112072468,-0.00677159244194969,-0.0127886107089016,-0.0136479120788762,-0.00586657635699306,-0.00231862303396591,-0.00540133971652934,-0.0047833851380209,-0.00431876724489622,-0.00697676784298473
"2789",0.000496894034754725,-0.000200421867491585,-0.00568721819137019,0.00869736012161448,0.00590119617495111,0.000290716960401394,0.0157743956196363,0.0108145514365519,0.00670346198651117,0.00117094409959151
"2790",-0.00113536131098901,0.00180508826730907,0.00492531702865096,-0.0135214025441646,-0.0144925001738412,-0.00515866512352137,-0.0166751166592216,-0.0116499679460911,0.00329028588656044,0.0099413840415421
"2791",-0.0217697732520364,-0.0248248302742261,-0.0147034489017981,-0.0256257087904905,-0.00927923413362441,-0.003703690603992,-0.0102264302527058,-0.0204474722144211,-0.0131178879376496,-0.0162129851678451
"2792",-0.0418226911338898,-0.0412646682717752,-0.0473364173446654,-0.0350662512799548,0.00944989378994521,0.00821754889795101,-0.0321737267006785,-0.0351179517259679,0.00253184589391431,-0.00941735710162106
"2793",0.0197025640752655,0.0220555811820418,0.0242547356410052,0.0325374142335042,-0.00621345010939733,-0.00436662637637231,0.00351351275606104,0.0132348638700877,-0.0104964249901067,-0.0059416896181449
"2794",-0.00542505657362713,-0.0121516439321309,-0.00888017478551673,-0.0315120922350867,-0.0095033108608189,-0.00292359192773639,-0.00390548543569169,-0.00979669282439399,-0.00470566289772678,-0.0113568727483593
"2795",-0.037508841823075,-0.0250264190866136,-0.0296996723611453,-0.0346504028044362,-0.0010938182066359,0.000880146914798541,-0.0294710905370531,-0.0228309091035417,0.00152257391199151,-0.0102780351854992
"2796",0.0150214684649379,0.00348049220847235,0.0100889318260831,0.0159773176338815,-0.00631906412200423,-0.0017581192847731,0.0207549932720998,0.00882635476948135,-0.00168031681036196,-0.0146611405460728
"2797",0.0146845487537146,0.0123563762224532,0.0194685184239136,0.0157259662919813,0.00440921234092895,-0.000293307855694813,0.00300209094459047,0.00823507924478606,0.00480889648494576,0.00619967137823907
"2798",0.00248748147186628,-0.00214141943161628,-0.0122883253488856,0.00763523333075766,0.00447393189712764,0.00166334090437292,0.00761898917788639,0.00306240770178601,0.00566322870710945,0.00184840363382421
"2799",0.0134960680770086,0.0199570598026457,0.0151311387441788,0.0250473335726789,-0.0110933936942155,-0.00605698474083893,-0.00486066339009539,0.00610725748548169,0.0170526171152821,0.0153751344041695
"2800",0.012760181040375,0.00736388263919796,0.00480281612409783,0.0205338436709566,0.00339931714313435,0.000294681310944789,0.00990475458700035,0.00354078218768983,0.00116984328690162,0.00181718054121949
"2801",0.000293001736948684,0.00104423205853443,0.0153289219798118,-0.00321930591981423,0.00542051023069767,0.00235836834315206,0.0084644294633518,0.00579614585769561,-0.00327158423151652,0.00181375993405042
"2802",-0.00626140829734767,-0.0110577048424919,-0.0081169163930529,-0.0137262658058962,-0.00438034452654379,-0.00107839108389263,-0.0123902463639525,-0.00501122720061853,-0.0134417084514044,0.00301758450131029
"2803",-0.00497401454988378,-0.00443038753556313,-0.00998359664175619,-0.000818733360381296,-0.0122686685780864,-0.00294380715821618,-0.0165925046468381,-0.00805832788470062,-0.00459437586492994,-0.00120347674362009
"2804",0.00129598820114318,0.00508574411912233,0.00462890258879578,0.000614547760000361,0.00299836535286691,0.00137784033983102,0.00932794522339764,0.00279237838048774,0.00509310026760779,0.00903620732628263
"2805",0.015939311217315,0.00674677877782326,0.0146452468928338,0.0178097270464288,0.00888196072361658,0.00383335898514003,0.0169884926047073,0.0151898180315773,-0.001266856660328,0.00656719708467035
"2806",0.0116122815866757,0.00649226721158258,0.0129744503559168,0.00925173527331835,0.000338497639371216,0.00117502735345032,0.00347442457240699,0.0107231299533774,0.00245757097239219,0.00533812706251435
"2807",-0.0124864662228336,-0.015813794587854,-0.0136086886540313,-0.0290953160990813,-0.00143848707725525,-0.00312962588857635,-0.0210412980298248,-0.0217121827869671,-0.0104389089072101,-0.0100296031652974
"2808",-0.0101301658331685,-0.0109936063534085,-0.00876479864484636,-0.0143678235145276,0.00635594360691427,0.00235458323756998,-0.00244856689470918,-0.0103403043620608,-0.00103889557353709,-0.0107270933030973
"2809",-0.0145405747944843,-0.0106882346236744,-0.0289831854364998,-0.00187409358412649,0.00682625361080791,0.00430326695042971,-0.00313677867036932,-0.0030580862187346,-0.00223999200000002,0.00180720426467462
"2810",0.00515507921978742,0.0010804266323452,0.011298488161092,0.00417270000809533,-0.00812946735835784,-0.0037092150868695,-0.00177832585496751,0.00996927463359421,0.00537201727572145,0
"2811",0.0115578786077724,0.00669106645000928,0.00450227112760815,0.00145442137021412,-0.00270365918772975,-0.00127349788860553,0.0112376747904404,0.00202489175458398,-0.00167476674116562,0.00601333289763395
"2812",0.00253499378666278,0.00578906262570289,0.00614206245825821,0.00933608786372431,0.000931826186480134,-0.0000980157578307495,0.00636929597579083,0.000252301787886822,0.0107844623741811,0.00358632258656688
"2813",-0.00036654415477666,0.00255796976865419,-0.0084143679383587,0.00102773104379228,-0.0011002914969469,0,0.00511694114217565,0.00505069551516635,-0.00640162812298772,-0.0107207044128849
"2814",0.00483926818293945,0.0017012067141311,0.00615642195838562,0.000205361237735291,0.0057622760728655,0.00206023272359324,0.00509124232469405,0.00427124564813286,-0.00238627901379029,-0.00602051145286409
"2815",0.0174022462160019,0.00466989256363326,0.00248039914419707,0.0213507737090066,-0.00657169094784615,-0.0021540572056542,0.00626508690748384,0.00150122073314418,0.000956809136609893,0.00969115162118062
"2816",-0.00125534272302419,0.00169015006004791,0.000989866878621681,0.00241206881283373,0.00576695607660338,0.00235476687815117,0.00503358239918494,-0.00299782292878914,0,-0.001799615516479
"2817",-0.00646244141989138,-0.00864790397901016,-0.00164796868411621,-0.00902345035104712,0.0050596544658037,0.00166399561032327,0.00158167380159968,-0.00375835384480216,0.00191172533127504,-0.00300482847068939
"2818",-0.00513159086909876,0.0025531404340795,0.00429179476726005,0.0016187407059256,0.00880937676022775,0.0019546916514972,0.000789710125046916,0.00653913328313815,-0.000636047071363111,0
"2819",-0.00108984773145981,0,0.00197238584226134,-0.00363622698246591,0,-0.000390267844034731,-0.000262914169474771,-0.000749421812443196,-0.00636431996096221,-0.000602764527766642
"2820",0.00108449169296088,0.00190998460182179,-0.00442922220812758,-0.00223040445306399,-0.00357638830737694,-0.00117072779446992,0.00591866066007696,-0.00248821650028264,-0.00240195352438821,0.00361883050760348
"2821",-0.0135304102107144,-0.00635447077065177,-0.0169714479616608,-0.0107700987092679,-0.00317163889586658,-0.000976727775955033,-0.00928341713327818,0.00428301152395894,0.00216697435259983,-0.0066105484132043
"2822",0.00170057771328791,-0.00127907682321704,0.0056990435460329,0.0110928673837922,-0.00401887698994263,-0.00195591993876698,-0.000791873253258912,-0.000501701837463342,-0.00448470398451106,0.00665453856253961
"2823",-0.00191910315295307,0,0.00133337923223076,0.00589176197106323,0.00109273645444574,0.000686018519886478,-0.00766092770013427,0.00175699999820145,0.0174563996051227,0.0180288471202825
"2824",-0.0249971997724318,-0.0217716249269214,-0.00915451881450002,-0.0333265052548793,0.00990952185740834,0.00411198350094355,-0.0057978002928083,-0.0122778111565018,-0.00395319408713168,-0.00767416064361603
"2825",-0.0213146096989234,-0.00654597624905073,-0.0209978325912273,-0.020267538678627,-0.000748718533341686,0.00136515392485292,-0.0159286125951645,-0.00659525167862529,0.0129385454928113,0.00892313813065582
"2826",0.0273590998538378,0.0197672304628045,0.0142416211546839,0.0324163631285819,-0.00382771857705311,-0.00272642202420836,0.0126199202637274,0.011491256102617,0.0052503565139852,0.00058967534721921
"2827",-0.0170116932557874,-0.0105535331088027,0.0023684852156145,-0.0181781036783262,0.0106926913831451,0.00566255660057191,0.00270935240357972,-0.00580659295975516,-0.00615841133581552,-0.00412480965262829
"2828",-0.00295502651916479,0.0065303024787573,0.0113079516645314,-0.00504954920778455,0.00264466443646572,-0.000193769447617398,0.0193190882587961,0.00761814909446001,-0.013804965311867,-0.00414207687878376
"2829",0.0127777591729423,0.00843426796134028,0.0126836140875812,0.0209346896059961,0.00486341724206119,0.00203891002917889,0.000265335979873216,0.00856829961814642,0.000477197157149556,0.00891265673453767
"2830",-0.0215845217024997,-0.0139395896698792,-0.0201053970957178,-0.0180198173174558,0.00197315381616914,0.00101951793576149,-0.0137806143793892,-0.00849550756393036,0.0116861514294764,-0.0135452839627221
"2831",0.0128168604912315,0.00587215939248975,0.0126134320955464,0.00991353298712161,-0.0077124369824576,-0.00320025897649878,0.00658339742385339,0.00579614173714349,-0.0075436035275247,0.00537306070353027
"2832",0.0106993116851064,0.00410798126170087,0.000996485773134381,0.000417756585292972,-0.00206730901748897,-0.00058379271038167,0.011211994517025,0.00927101828038945,0.00118760092190962,-0.00415671294288755
"2833",0.00789207674650649,0.00969003753246334,0.00497759029041855,0.00250513957860665,-0.00745700547070871,-0.00253110665672929,0.000924140000308604,-0.00099302847527305,-0.0051403243607826,0.00477048083169485
"2834",-0.0222861478379862,-0.00447857506778382,-0.0156843078659947,-0.019575048211695,0.0109357368293028,0.00439179243795396,-0.00896760497511584,-0.0042245880270646,0.0046899521934034,-0.00712168600849572
"2835",0.00492854259266684,0.00921174886719456,0.00888969084967051,0.00106200325364436,0.00165172857803375,0.000194528346282308,-0.00172976097264299,0.0069876874082706,0.00340217583196578,0.0125522520913601
"2836",0.0159000913215626,0.0123114974887999,0.00548620802676125,0.0195204076652649,-0.00181371384458029,-0.00174881558476025,-0.00386547698528561,0.00669120463516437,0.00236558113862162,0.0171191926377148
"2837",-0.00524196958706014,-0.00671001887924771,-0.00248011030209383,0.000416168520056992,0.00355111783171225,0.00097323793608628,0.00227451354646058,-0.00147682941372496,0.00778790101192817,0.00754505613080703
"2838",0.00822695834483378,0.00654434805393977,-0.00165754657118689,-0.000415995395868785,-0.00732420549428514,-0.00359724472581213,-0.00947912179075727,-0.000246796703604613,-0.0116306142250363,-0.00403226212851959
"2839",-0.00293323411855484,0.00167765284905874,0,-0.00998954109458905,0.00232125396807614,0.000878242135959217,0.00350450575872396,-0.000739703868756214,0.00655499905492807,0.000578361080894707
"2840",0.00822186394938385,0.000628235458893345,0.00282255446628543,0.00126130348432207,0.00033083974665038,-0.000487278620449172,0.00483538522000648,-0.000493529945614246,0.00141231858954072,-0.0034682796207488
"2841",0.0106983560178859,0.00732372902915546,0.00380794384236816,0.00209947993032578,0.00272843789526611,0.000584956013209625,0.0129663193790202,0.00691361400480672,0.000940241344673742,0.000580157907066337
"2842",0.000740512382854996,0.00332367002692657,0.00676229852292543,0.00858992658884405,-0.00799856149361833,-0.00389878954899159,-0.00171560881456234,0.00294264554497636,0.0007827632093933,0.0185506490623992
"2843",-0.00554759753740641,-0.00434781162536779,-0.00376801795121773,-0.00581627965610532,-0.00814642255978359,-0.00274008095444689,-0.0142765673457621,-0.00537893545418178,-0.00195541653430453,-0.00398412652387103
"2844",-0.00847919249608164,-0.002703380596774,-0.00197349631796861,-0.0125366965807603,-0.0072074042570357,-0.00333645366387325,-0.0085822859303768,-0.00147522824371837,-0.00760188883388535,-0.00171426242459438
"2845",-0.000150213093432328,-0.0012509839035052,-0.00131808209186812,-0.00804049847192467,0.000253187247631237,-0.000984640495977351,0.000676224092121425,-0.00664673000454929,-0.00797594585744166,-0.000572402055533772
"2846",-0.0134674082783902,-0.00501038337509274,-0.00362970807123142,-0.00469291663635385,-0.00455720606142107,-0.0011822165403933,0.00243332354726267,-0.0014869440669274,0.0048559145473035,-0.00515456898568611
"2847",0.00247179469546688,-0.00356704010869913,0.00314620767400786,-0.00771532453309653,-0.00669778401011123,-0.00217102440833949,-0.00215746544689832,-0.00297863741849524,-0.00649607051027323,0.00172709207715172
"2848",0.0101655796080096,0.00568535665343961,0.00610757333710432,0.0144708240500335,0.00699888030785201,0.0028675908634157,0.0121619072212578,0.00896181910658189,-0.00350851595539381,0.00517234311863457
"2849",0.000938887213706607,0.0012564934934467,-0.00278914325012358,0.00617406268653053,0.00771323753248687,0.0016762095145697,0.0129507258846007,0.00542827345013741,0.00424100980842601,-0.000571629824671294
"2850",-0.00769060834566704,-0.00460066977743145,-0.00230333961543439,-0.00719406896961605,0.00176631806113092,0.00108287069809498,-0.00303152545045682,0.00147255019543868,-0.00725102788844623,0.00457659625192264
"2851",0.00177684561061509,-0.00546214739421425,-0.000824562303778476,-0.00490213524114247,-0.00360149257951248,-0.00156627700012657,0.00700677831788399,-0.00196040777034256,-0.0070631433361632,-0.00569480027258995
"2852",-0.00671747956733915,0.000422425488944889,-0.00594158921476218,-0.00792447893320547,-0.00109778271648753,0.000197408226883411,-0.00341329485630337,-0.00785665916398792,-0.000484981007881191,0
"2853",-0.0022036630441431,0.00358945340659989,0.000996154859596698,-0.00215887925767,0.00448069575086829,0.00256465456414601,0.000395271245605011,0.00470168945845573,0.0050950019394258,0.00630014665445522
"2854",0.0129463844822892,0.00189366769066335,0.00729812011356712,0.00454354902206533,0.00151504985586604,0.0000985917880074183,0.0105345628748217,-0.00123155292522592,0.00209206631873249,0.00682990607890632
"2855",0.00338333640514321,0.000839973919101844,0.00115261794462995,-0.00581533917364363,-0.00159652212568206,-0.000492117568264616,0.00547309892696357,-0.000739703868756214,0.000240878430697755,-0.000565341543789177
"2856",0,-0.00125894867865139,0.00312497431957759,0.00563262497616468,-0.000925903540612394,-0.00167347554345687,-0.00492502723982557,0.000740251435606964,0.000160520189451674,0.00282807382389816
"2857",0.0096657310203867,0.00693275341763067,-0.00852590449053758,0.00193868949711362,-0.00598233994507213,-0.00226771503792544,0.00612158313394118,-0.00271256615687376,-0.00208679676015089,0.00902412904987493
"2858",0.00935065368784427,0.00479862323420055,0.00578786881296245,0.0208557366628574,0.00805239546099479,0.00207537638205069,0.00919085645063378,0.00642936562616536,0.0068366282178618,0.00503079018948172
"2859",0.00305109719263497,0.00145357320627082,0.00756331315941106,-0.00168479236897423,0.00252242280336334,0.000098897971329448,-0.00410480328970808,0.00147424365141879,-0.00143792938169041,-0.00611782543922279
"2860",0.000476699200071318,0.000414719796316687,0.00554831503593278,0.00126573791893736,-0.00528396413902366,-0.00216976150176318,-0.007341486425679,0.00318932918786641,-0.00408001599999996,0.0072746624522757
"2861",-0.00688720460594672,-0.00518143503062052,-0.0102239366373938,-0.0206489738617461,-0.0113828206732643,-0.00553404056059192,-0.0147917615729904,-0.0124724996585887,-0.0161458352662196,0.00111115316920229
"2862",0.00420521429671328,-0.000833391568088149,0.00295134516227358,0.0150603626756978,-0.00383778065308749,-0.00208709189831713,-0.0028972936930739,-0.00470506601162779,-0.0015512899685346,0.00554942804543024
"2863",-0.000844882788980539,0.00291908983676348,-0.00016354853325351,-0.0152608456836426,-0.0050513025978639,-0.0005971571841632,-0.0051511279010189,-0.00497661086127921,0.000572409840768451,0.00110373765033045
"2864",-0.00249995111001211,-0.0037421853060261,-0.0024526038430468,-0.00839421111776262,0.00860501286297621,0.00388589509742188,0.00225692683542178,-0.00300074809421613,0.000408654785807094,0.000551146903571942
"2865",0.00751865345251845,0.00605172049521308,0.00114744814943202,0.00607768299256706,0.000511889428863155,0.000694737126592404,0.010729620934834,0.00652116476626596,0.000571840517217925,0.00771362090786609
"2866",-0.00278015793974573,0.000414981357037991,-0.00229214625070806,0.00345189365426868,-0.00153481072094808,-0.000396736305964929,0.00131076555007614,-0.00249207039241228,-0.000571513702526616,0.00109347875985599
"2867",0.00275115315161978,-0.0143065028113245,-0.00393831564472891,-0.000429948382092094,0.00725945015133567,0.00456446004717481,0.00850805076542471,0.00174886611267899,0.00106198019567105,0.00546159048228656
"2868",-0.0020484537710953,-0.00294478814796262,-0.00609549948205823,-0.00537736026530367,0.00796986337984529,0.00256811340093832,-0.0024659658871018,0.0017455199979941,0.00856858977828789,-0.00651827470529265
"2869",-0.00238275568404434,-0.00886086605959002,-0.00331502383898108,0.00410901044808032,0.00622506778967957,0.00394088665887682,0.00338255320695846,-0.000995660208102045,-0.00307465824337438,-0.0147621883463144
"2870",-0.011501018414054,-0.0266069700277557,-0.00665242983255987,-0.0232609694866488,0.0219025584633226,0.0107946093006976,0.00298240340720324,-0.00971831350350905,-0.00016230013929297,-0.0094340048311472
"2871",0.0133447008827769,0.0177126656087776,0.00703177145575529,0.00793828594577373,-0.00670832443586078,-0.00427144959837289,0.012669937810956,0.0103171095682877,0.00146116565531007,0.0128852670219088
"2872",-0.00612585884407868,-0.00429740051206096,-0.00681627947394037,-0.000437588819436785,-0.00164706639835122,-0.000487713306080884,-0.00178743045535878,-0.00423426240402824,-0.00218857901786706,-0.00276550571138057
"2873",0.0098177613354451,0.00820028466320899,0.00686306000900805,0.0140076530788793,-0.00528355459636565,-0.00369449122812138,0.00345313941450187,-0.0002500538904181,-0.00495532095784434,-0.00665559702864238
"2874",0.00475134660460008,0.0025683723853327,0.00598498264724134,0.0101443746153518,-0.00723175897656358,-0.0035319247971668,0.00879427713777425,0.00850625094186741,-0.000979631006280179,-0.011725247698573
"2875",0.000727706387750882,-0.00170792321591939,-0.00181781010645554,-0.00769226736559092,0.0023441446780379,0.00255973305128387,-0.00126356772686764,-0.000992085578002566,0.00392248907601966,0.00169489199511852
"2876",0.008360517033281,0.0100513193610465,0.00430458476687834,0.0150732431789955,-0.00810307244855712,-0.004026322758102,0.00113853331196623,0.00645603936440908,0.000569800579077073,0.00338416449252255
"2877",-0.00010836279468851,-0.00804569104553687,0,-0.0152736166661149,0.00968540703412835,0.00423988444160606,0.000631911653399708,-0.00764853820446454,-0.000488097957827893,0.00393474064972654
"2878",0.00295635272570571,0.00128071495603455,0.00296733200144605,-0.0019386894971134,-0.00300293544153052,-0.00137465086020516,0.00290422520146993,0.00198916608174371,0.00122090996890023,-0.000560017988806005
"2879",0.0013301492527138,0.0100191784524664,0.0031229199110463,0,-0.0018405143636524,-0.000983190814357493,0.000251868087530971,-0.00198521715511379,0.00178848058225367,-0.000560216466350849
"2880",0.00129240802321462,-0.00654287527411035,-0.00622639528827296,-0.00259021433295448,0.000251262202932256,-0.000590418996850861,0.00503527568331963,-0.00447522211833762,-0.00332713616829172,-0.000560415101785283
"2881",-0.00319104591193275,0.00212442623563658,0.000824357453331759,-0.006708550567047,-0.000502600759204608,-0.00118184413266031,-0.0201652223218267,-0.00174825287656166,0.00301255495847585,0.00392579808687055
"2882",0.00251778626473875,-0.000635933354659834,-0.000988372808864546,-0.00675383613288982,0.00829989825987454,0.00315497021691402,0.00997047556798836,-0.00375289260492317,0.00154229236882375,-0.0111730327424138
"2883",-0.00127577189903405,-0.00615187749336843,-0.00527710566289485,-0.00789649618266186,0.000914529354048232,0.00078624139252037,0.00101241255249085,-0.000785564839732911,-0.0165342928319248,-0.0242939171124082
"2884",-0.00205663427956704,-0.00917829992149188,-0.00729435175196147,-0.0121600435377336,-0.000913693754289291,0.000490867379582705,-0.000884929103836085,-0.00532588341018669,-0.00189545910319633,0.00868564270287542
"2885",-0.00383284486426139,-0.00844302447930101,-0.0106025263375158,-0.0110385365329475,0.00582012714297719,0.00265033672347803,-0.000126571512946039,-0.00535443000142866,-0.0025596399755623,-0.0103329868542164
"2886",0.00170603388159174,-0.000222327869539907,0.000340229790960933,0.00432799167314668,-0.00876230618779028,-0.00323055726918631,0.00974577416649436,0.00281974159281484,-0.00447020684262733,-0.00116019641551013
"2887",-0.00626892992557282,-0.00778280754177485,-0.00374091970909207,-0.014062025855378,0.00525365337958816,0.00265182631369498,0.0051390730058396,-0.00460111609617586,-0.0017462081864924,-0.0075492592332711
"2888",0.00182322236409749,0.0136708275846726,0.00494967657681289,0.0103517866246738,-0.0000828965372120516,0.000195754812141402,0.00635976226071966,0.00950181667543837,0.00241560177220479,0.0198948260359761
"2889",-0.0136129250202861,-0.0148129573751133,-0.0135869449850791,-0.0134333296923523,0.00224004036016368,0.00137130425035581,-0.00346937890700683,-0.00661430791144613,-0.00373938021403952,-0.0114746066791805
"2890",0.00221405145246645,-0.000224517956754711,0.00585391533729251,-0.00392353291190339,0.00140737402520563,0.000488769306627779,0.00395490136323895,0.00409734190998479,-0.00525479193639833,0.00986655672432346
"2891",-0.00828419620646703,-0.00965215931303987,-0.00667580805012269,-0.0192307060310637,0.00942399006010897,0.00381255341324604,-0.00537780435158819,-0.0119865883777778,-0.00570182784333684,0.00517234311863457
"2892",0.00571758137050637,0.00249327699313673,0.00120625694266696,0.00850463797393841,0.000245698682666218,-0.000974112888210366,0.0106877861331427,0.00309749861242348,-0.0030359334957677,-0.000571629824671294
"2893",0.00143964913367833,0.0108522903964099,-0.00327014050228458,0.0149918615587585,-0.00343875588480536,-0.000779803803281132,0.002488278930314,0.00720533848771754,0.00363729484319664,0.011441608389076
"2894",0.00213798971085666,-0.0071571726665195,-0.015886730748347,-0.00992393790329249,-0.000782335060692363,-0.000683878380211667,-0.0059568523859741,-0.00715379298776975,-0.0100295236404632,-0.020927723011414
"2895",-0.00353136784413066,0.00585716477268994,-0.00122834243369629,0.000699393080512367,0.00535642938978387,0.00254259499106446,0.00749040866222939,0.00591879927639893,0.0101311340893167,-0.00115526692314427
"2896",0.0081579629061912,0.0132139607747448,-0.00158109653987959,-0.0025624776781743,0.00286870827895225,0.0000975245433632033,0.0130112607724606,0.00690711884110784,0.0033712683797511,0.00578367033561245
"2897",0.00845823997811235,0.00486272931530385,0.00651063894172665,0.0137786872673766,0.00326937941640981,0.000877726814959345,0.0041589385658245,0.00685982653826867,-0.00159598484008439,0.00460028213185626
"2898",0.00900450912316164,0.00637940796327596,0.0138112131044292,0.0179682602027407,-0.00643590599488719,-0.00253367541016158,-0.00889254501115855,0.00454181517932439,0.00243985358876109,0.00515173632649257
"2899",0.00359830727478805,0.00240435316504195,-0.00379381778606458,-0.00226304026398017,-0.0000820042372181584,-0.000781344691433317,0.00307289041058634,-0.00276307776301643,-0.00184642884017738,-0.00227787321992068
"2900",-0.00731444891761168,-0.0183165802365851,-0.0138480069567707,-0.0195054890978937,0.00385409382883162,0.00205323885430309,-0.00306347668246576,-0.0130981942351691,-0.0108467249642648,-0.0348174624831071
"2901",0.00906587724015617,0.00888490797179586,0.00105318776646834,0.0136479093322253,-0.0000816361281665845,-0.00039037506951034,0.00294993157210843,0.00535989641536494,0.00416523294938154,0.00532240485517366
"2902",0.000787469804602203,0.00286217023764235,0.00929340731441486,0.000684613418322266,0.00253239168608554,0.00165923314991701,-0.00343122337328017,0.000507484532478397,-0.00440189632782273,0.00176480282097224
"2903",-0.000893995645425583,0.000438998876224783,0.000347482137547761,-0.00547316034756373,-0.00415552949653897,-0.00165648465566393,-0.00455018446169964,-0.00050722712255924,-0.00051014369092639,-0.0211392979429703
"2904",0.00404512475811125,-0.00175531745046498,0.00885713115842157,0.00733769954945762,-0.00188205838403299,-0.000585709871796181,-0.0053117445137002,0.00025375704189079,-0.0108039469807585,0.00119974367765274
"2905",0.00210384043731926,0.00241800239180567,-0.0015492514195341,-0.0011380616545571,-0.00401740168164133,-0.00078151278318972,-0.00471932813855147,-0.000761432522448424,0.000257989338303899,0.00898741846514817
"2906",-0.00377170444516062,-0.0035088794364313,0.000172324678149316,-0.0123062861600025,0.0063382627354609,0.00273727103648369,0.0101071368465722,-0.00558788648981534,-0.00429885657809059,-0.00118763226939633
"2907",-0.00114275174950984,0.00572191416465584,0.00310299052674368,0.0143053676662157,-0.0122689233543702,-0.00350962521972509,-0.00840019876362497,0.0109835278004751,0.00647612479882786,0.00713438888152895
"2908",0.00185920762884018,-0.0026258088643184,0.00498362949030384,-0.00659694135726008,-0.01233855257828,-0.00489145808644642,-0.00249158193214305,-0.00480053252263646,-0.00480437551139967,0.00354192497063477
"2909",0.00503224530573521,0.00680104410095805,0.00410399232954206,0.0146555262513359,0.00343759871950722,0.000688137698376501,-0.00487088526103863,0.00330026000714256,0.000344836206896515,0.00529404521019172
"2910",0.00852252909881135,0.00740915819619281,0.00647136586295316,0.0162489511684716,-0.00158762269826906,-0.000687664490516604,0.00815805310920714,0.00607284575531408,0.00551533087284284,0.0134581601662647
"2911",-0.00235915988975033,-0.00605658559781785,0.00253814585636225,-0.0111036366250894,-0.00192476033885136,-0.00108127578921469,0.00273848404298027,-0.00829974511461873,-0.00779913438464175,0
"2912",-0.00677645897444556,0.00195861894376503,0.00303797994868105,0.00359306258122016,0.00167674039402033,0.00157447001563349,-0.00968342566988656,0.00152188340629,0.000518312184114356,-0.00404145601756001
"2913",-0.00522344595697533,0.00260641752044988,-0.00757203371578696,-0.00156634134081779,-0.00343179837588425,-0.00127721197124575,0.00137886137094734,0.00177244940209786,-0.001554001527169,0.0057971412257396
"2914",0.0049293880517407,0.00411594729160569,-0.00762964859415105,0.00537880538566227,0.00545971014359981,0.00137736873617378,0.017150650417022,0.0045500875373321,0.002939870247473,-0.00576372808007275
"2915",-0.00167044988110077,-0.00755108687589467,0.00649237312385487,-0.00891663630124695,-0.00814673819296985,-0.00236273309191115,0.00332319600231057,-0.00603957740415628,-0.00732820945474966,-0.0144927933996526
"2916",0.00544752384737146,-0.00913041704563189,-0.0056017226437195,-0.0132703596597438,0.00143493917259119,0.00118415927709714,-0.00331218894923557,-0.00278452741053248,-0.00538476641814112,0.00588239354001052
"2917",0.00428470364865308,0.00197451829983053,-0.000170742437803573,0.00775021287010258,0.00497364919049725,0.00256259771018286,0.011815689250541,0.00406197440236533,0.00349284850225762,0.00350872377936784
"2918",0.00366712895856969,-0.00459834560517824,-0.00751230324076779,-0.00769060901315,0.000587229067717798,0.000491620391037006,-0.000608215780008359,-0.00455135561179631,-0.00513397154775463,0.00174822784108608
"2919",0.00330250063363713,0.007919177941347,0.00842932548427022,0.0102574973229728,-0.00519771071736319,-0.00206348434415349,-0.00352970183947898,0.00330184825861335,0.00227406625952842,0.00756249299486456
"2920",-0.00042027250947807,-0.00174583209606982,-0.00102354326451159,-0.00135368509011013,0.00101144001263043,0.000886310762925113,-0.00598528929470088,-0.000759151345356535,0.00279263470783264,-0.0121246057469363
"2921",-0.00136605935674672,-0.00349811625098051,-0.00375681954293638,-0.00293714998956685,0.00841820052000508,0.00275459079786922,0.00122885146199159,-0.00354713776473559,-0.00147947083876176,-0.00409111864171874
"2922",-0.00670023283016929,-0.0223781360547248,-0.0143983264793029,-0.0213008246955886,0.00726270051630706,0.00431642662645326,-0.00895911748446021,-0.0142383190530269,-0.000435732969073177,0
"2923",-0.00374339377099975,-0.00269317506082445,-0.00591303567916779,-0.0164388521620874,-0.00207196835831902,-0.000293018002287759,-0.000495444462781491,-0.00464313259048665,-0.0150841657496876,-0.00528167780563416
"2924",0.00638067780056994,-0.00180014049460664,0.00402367277510551,0.00612056864552768,-0.00224235839321385,-0.000977060399296126,0.0054516872629895,-0.00259117229589978,0.000973804895306296,0.00176976566726261
"2925",-0.00746727626039767,-0.0171326500713145,-0.0121971790251788,-0.0287788217740838,0.00582646898447581,0.00244507047860476,0.007516977970077,-0.00545586132431675,-0.0166268506235074,-0.0217903474683254
"2926",0.00809122419556307,0.00711028648350065,0.00546832797570018,0.00626359403128696,-0.0000826489479700543,-0.000292756147620254,0.0080722612496682,0.0070532728526429,-0.000809461267929579,0.00782656574689478
"2927",0.00352050069591581,0.00592109566641352,0.00333332108057283,0.0105338086742019,0.00124127433318066,0.000390537073468034,0.00897851127177263,0.00648493752049695,0.00927091825870252,0.00418166710267975
"2928",0.00214017420440227,0.0070183390163181,0.00402165305989932,0.00450144991626389,0.00669545906463953,0.00312205171942459,0.00156333726958824,0.00670124983994635,0.00499424788176883,0.00178462762613107
"2929",0.00234500098897206,0.0107913902540804,-0.000174137600244095,0.0127357463835172,-0.00336683131987436,-0.00136158768085326,-0.00672349889321777,0.00179196195203257,0.00292834319055202,0.00178144840409455
"2930",-0.000593669041566547,0.00333630753827485,0.00418053618825653,0.0079180681504154,0.00395471726013552,0.00185038701406204,-0.00556041908456295,0.00178887555896212,0.00221199793519733,0.0142265489565536
"2931",-0.00132781620327982,-0.00753724582125226,-0.00416313206400643,-0.0161736309637286,0.00155921267539982,-0.0000971439742371016,-0.00218812617711261,-0.00612245007041168,-0.00944645562231283,-0.00175333656073662
"2932",0.00601839755824862,0.00826450540633195,0.00348373800005097,0.0185532675687157,0.00196641331622982,0.000291389432164557,0.00511662374559818,0.00487692830272146,0.0174688685597737,0.00761113664734459
"2933",0.00789538276587964,0.01329215570008,0.0151015177748783,0.0142954724031088,-0.00572411048929511,-0.00223528310872689,-0.00181803914636569,0.00791823002423153,0.00376657309857831,0.00348629761126173
"2934",0.000483135669854029,-0.00174913875113236,-0.00307798094467682,-0.00363707373761624,-0.00600386930136076,-0.00224029079289467,0.0106848453883506,0.0012671834674105,-0.00794132150942739,-0.00405309730294123
"2935",0.0053807283358025,0.00459914503374859,0.0036020648557773,0.00616004259249459,0.00132399142508288,-0.000292693952251954,-0.000961041943808638,0.00556808538852449,0.00457421710063333,0.0110464194354272
"2936",-0.00404820027983932,-0.00981024479372139,-0.00700737956938324,-0.0260770885376408,0.00214853860118192,0.00185514149854615,-0.0034873474907523,-0.0113264440264668,-0.00490366037400147,-0.00172510579944607
"2937",0.0000343615379649886,-0.0112286692586784,0.00206547968353754,0.0051222025042672,-0.0023088289085611,0.000195132628983741,0.00374079430326302,-0.0015274580468374,-0.00114393700408255,0.0011520579548232
"2938",-0.00172229852041716,-0.00823864841438737,-0.0123668525970063,-0.0194578998835503,-0.00578156403571373,-0.00228516454975392,-0.0105793195501543,-0.0114736089779459,-0.00510969949590867,-0.00575372044135014
"2939",-0.00269144130148524,-0.00583741609676891,-0.0106087140236498,-0.0144104766099495,-0.00266602303828112,-0.0000978570853215066,0.00461716616033758,-0.00438510738820364,0.00345346674931357,-0.00405098955429095
"2940",-0.00301008704104744,-0.00496834528193635,0.0022850973862043,0.000958672663338378,0.00367554597339481,0.00205544383740808,0.00387026956121672,-0.00103613396190749,0.00194141369572898,-0.00581049601876982
"2941",-0.00194329138106508,-0.00817061615771908,-0.00613824433627597,-0.00502869539834538,-0.00848924841423482,-0.00449339282829708,-0.0121686009780555,-0.00674280712148367,-0.00273029766839628,0.00233778208098223
"2942",0.00173841842630584,0.00892444495881795,0.0022939685604848,-0.00986766801977523,0.00369344034120611,0.000588834070536448,0.00634227098162965,0.00104446257042579,-0.000706535351765347,0.00349849440394534
"2943",0.00329745872558185,0.000453535916852044,0.0021126799143476,0.0021876344142866,-0.00761058834107564,-0.00362870955748051,-0.00206051626485348,0.00365159229875123,0.000618638963877371,0.00987802264203652
"2944",0.000242232140178489,0.0038540242942815,0.00193257686099058,0.00509326148926514,0.00235953588913329,0.00118116957525394,0.000850246445169178,0.00545727852820677,0.00839071711366635,0.00690439346752192
"2945",0.00591446602666079,0.0072267467798881,0.00771521497057459,0.0135137029832089,0.00151326258970141,-0.0000985145725520553,0.00594596646588652,0.00361852911468374,-0.00359110105266014,-0.0108571717928199
"2946",0.000171932689684295,-0.00224212682878888,0.011310233141907,-0.000952381619472531,-0.00478504685348513,-0.00186802073115788,-0.00808202069411956,-0.00309043932730046,-0.00650496648198018,-0.00635450319835917
"2947",-0.00529438460150033,0.00269671196340249,0.000516245759894396,-0.00905626291129369,0,0.000197182097129822,0.00352648846863413,0.00258313929893594,0.00522035051903247,-0.00116289437072703
"2948",0.00542621113078434,0.00515448994376211,0.0239036677702777,0.00961991547343199,-0.0104597769855843,-0.00413628551263578,-0.0035140960494382,0.00669973388760292,-0.00149633833732643,0.00931320734642194
"2949",0.00106571325221916,0.0022297229707231,0.00352706433311556,0.0138162017417283,-0.00596692967861345,-0.0016811115266796,-0.0132556784519243,-0.00358357233548057,0.00387865825319711,0.0063436269774495
"2950",0.00810384392973007,0.0180199891534922,0.00267781160323333,0.0110432348170457,0.00463084684067505,0.0000988751366655105,0.00998277212183019,0.00796306787491363,0.00342465762446409,0
"2951",-0.000913703954341205,0.000437053336256543,0.0021698907544121,0.00464789895819173,-0.000426880409003849,0.000396088802794958,-0.000487980376124297,-0.00790015837753066,-0.00682592999455489,0.00229223237918608
"2952",-0.00332199113806719,-0.00480553247648829,-0.00449701007835257,-0.0113346384510487,-0.00256178780825966,-0.00108896971833317,-0.0175803204703652,-0.00363341751416846,-0.000176200549408811,0.0148657296621684
"2953",-0.000927725817140512,0.00570672717900034,0.00752894363583967,0.00397739984552636,-0.00102750429768617,-0.000991078829118863,-0.00161558419687635,0.000520875315407565,0.00158633117488027,0.00225360625707682
"2954",-0.0029921110305271,-0.00152767207110382,0.00481558080486466,0.00209739648256679,0.00702777934771914,0.00327412718392162,-0.009150392858292,0.00364488888474312,-0.00527935758417319,-0.00449707787132436
"2955",0.00279391060732648,-0.0028415941282719,-0.00264416156410996,0.00488368210831314,0.000680785811689288,0,0.00266395575699319,-0.00181584090100562,-0.00884564328582993,0.0045173929391471
"2956",0.000103355039405617,-0.0120560934421382,-0.00198842173542801,-0.0067114454611289,-0.00263654999424046,0.00049464328797022,0.012398401104794,-0.00597714951804718,0.00633644784462883,0.0101179045278676
"2957",0.00347433004632824,-0.000443767781570736,0.00680728566917077,0.000233193775287965,-0.00734136243785566,-0.00253557419160599,-0.0082476746575314,-0.00261436105271873,-0.0016850123858636,0.018920451388869
"2958",-0.000583014337249277,-0.00532729692142153,-0.00230872829635054,-0.0125787105540468,0.00611301702997924,0.00258173631688763,-0.00138596604495567,-0.00996076362965514,0.0115483965532557,0.0032769655314917
"2959",0.000548971097974249,0.00379362991845111,-0.00876031190949189,-0.00825661493485652,-0.0173711902300896,-0.00742805393761525,-0.00694013129167803,-0.00529514115536756,-0.00395191875071776,0.00925425988695894
"2960",-0.00781586789169908,-0.0131168523752082,-0.0135067253172619,-0.024976287464706,-0.00705402686830914,-0.00259428678097728,-0.0100382239260098,-0.0188980492309569,0.000529051323030272,-0.0107876155675189
"2961",-0.0055969743239298,-0.00698355539477002,0.000168998358354155,-0.00365940001988052,-0.00859490024491782,-0.00240101323706099,-0.00128346211674557,-0.00189912698355899,0.00281988008054612,-0.00218110757682066
"2962",0,-0.00930134053877563,0.00439416148064864,0.00146921334429262,-0.00336169506941386,0.000401234178543097,0.0132373102998853,0.0046209770739527,-0.0110720735218258,-0.00273220340393854
"2963",-0.00145931110281095,-0.00114498596158663,-0.0057210785661721,-0.00366755489746728,0.01011881588708,0.00190442278514058,0.00215630282740609,0.00865769857118615,0.000533117109177805,0.00712324725195068
"2964",-0.0316630856611556,-0.0194863491083777,-0.0245388303342789,-0.0296931006555894,-0.00272400454465194,0.000500461189002488,-0.0150614138955791,-0.0179719206779069,0.00248666967116651,-0.0195864096426023
"2965",-0.022026642799408,-0.0126257388721943,-0.0180430218303286,-0.0101164770643761,0.0121596861638875,0.00409988035228315,-0.0272422833805888,-0.00409721295427967,0.0256910176920009,-0.0149833186461571
"2966",0.0138884315388259,0.00189452091208664,0.00229680554504119,0.0293818029930653,-0.00348208604223921,-0.00119512123536181,-0.00198155873691475,-0.00191989894683298,-0.00475035416091174,0.00788721601174891
"2967",-0.00561684862075784,0.00165440619349044,-0.00299661960392028,-0.0106727545153544,-0.00043708540671783,0.000598234300082101,0.00542672032552827,-0.0010990055035438,0.00668226138985695,0.00223597067338011
"2968",0.0218655455761432,0.016045174304987,0.0185643341023374,0.025087932930921,0.00227231383174864,-0.0000997407617919777,0.0217220807927072,0.01980734992445,-0.0017241120689655,0.00446184972113572
"2969",0.000178544031832706,-0.00952147465525288,-0.000694307135204575,-0.0122370048470666,-0.00592939753014099,-0.00289003390326203,-0.00489630952254749,0.00161848590733493,-0.0000863730547572272,-0.0088840601011867
"2970",-0.0144410802707613,-0.0164127439990365,-0.0180649602538696,-0.026263634848785,-0.000350693287713422,0.00179918407104895,-0.00116534844222238,-0.00430921592047417,0.00112269625077555,-0.0112045023045214
"2971",-0.000542578628127455,0.00786644798719394,0.00212277041171594,0.00941469217474333,-0.00219395492915342,-0.00119727775758416,0.0076485846850296,0.00405731559710931,0.000776432035480168,0.00566582033804575
"2972",-0.00448882589582555,-0.00591294382871588,-0.00617833521058575,0.0108394278955557,-0.00131917758642075,0.000199483588825933,-0.0131225427176426,-0.00484919747850288,-0.00258600978215662,0.00112674514453537
"2973",-0.00509060926429417,-0.00713765240058739,-0.0115452033772638,-0.0109724731172089,0.00317013855455639,0.00259670201788764,0.00638780883763057,-0.00378981004948209,0.00587676091847511,-0.0219470914597191
"2974",-0.0302986858088858,-0.0282770272206634,-0.0319857724789125,-0.0322743826801382,0.00754928860205939,0.00537909725282937,0.00725379172475993,-0.0138587867377079,0.00231982990222379,-0.00690445268593698
"2975",0.0179405220730362,0.0128236259356773,0.0148506516774405,0.0192808225881316,-0.00418192652416227,-0.00237761995378172,0.012345823973527,0.00909341501222682,-0.0022287158502069,0.00405556430793319
"2976",-0.0175873876465605,-0.00413919628183257,-0.012804044255541,-0.0115029766548891,0.00603637903334042,0.00446900952608598,-0.0235008825501819,0.00191163642766612,0.00317865114813309,0.0075013995081854
"2977",-0.00554016390404155,0.000244403219094691,-0.00926438373853578,-0.0173261805948635,-0.00226077865176577,-0.0000990436483830903,0.0115777054478108,-0.0032708742507922,-0.003939359525718,-0.0103091969184586
"2978",0.0148182625301221,0.00855542226739647,0.0157097124036372,0.0194739635692553,-0.00496816099100028,-0.00217513895482979,0.0150464507810901,0.00464896563727879,-0.00438479072108655,-0.0052083811063095
"2979",0.0106810251323297,0.00799807654321216,0.00975869448882727,0.0108413375207497,-0.0050806176772209,-0.00247759622889299,-0.0103888809647954,-0.00816558587094796,-0.00561313456960799,-0.0133799887343048
"2980",0.0106418857262089,0.0158692551065303,-0.00237051789324716,0.0357507929454157,0.000926716471088218,0.000856082125329394,0.00371276069960258,0.0148187763431475,0.0128527570498871,-0.00707537594761776
"2981",-0.00592295702313017,0,0.00566630736485907,0.00641019629952,-0.0124327810820419,-0.00557047120757681,-0.00854601131046051,-0.00459704770842029,0.000171525340946443,-0.00237526453879289
"2982",0.00551682244645146,0.00070988138933159,-0.0036351424362201,0.00269475315255496,0.00392859498732312,0.000600050932030083,0.0146661680007374,-0.00135831710394774,-0.00240033429232178,-0.000595229963322619
"2983",0.00632788801721329,0.00165568009520234,0.0113097997830314,-0.00171012924285063,-0.000622514487150228,-0.00109953702926036,0.00431095121820912,0.00788895490527697,-0.00283579953160262,-0.00416921391002356
"2984",0.0214089823568411,0.0129870637160809,0.0104617605427528,0.0188447781534862,0.00133478393572894,0,0.012624471853111,0.0156546927075201,-0.0000861944149759264,-0.00239218884047798
"2985",-0.0018151997994994,-0.0114219425151936,-0.0064262878715009,-0.0259430255095329,-0.0000887130419781057,-0.00140116095217468,0.000373951426738017,-0.0087697203976933,-0.00215461520429727,-0.00599530645430091
"2986",-0.00976806956981913,-0.00377258736904851,-0.0100610660759985,-0.0184956434139217,0.00746583940042433,0.00390854574775346,0.00137116311004659,-0.00482576550211766,-0.0112281569461752,-0.0108564294470516
"2987",-0.0186852230533014,-0.0201183353447262,-0.0136115831132652,-0.0140702323940868,0.00652857731684442,0.00299512137295466,-0.00112029574983286,-0.00592668311857114,-0.00716281427770404,-0.00243899102184708
"2988",-0.00187094154879808,0.00748774456220058,-0.00367989743570774,0.0114679055068083,-0.000613720981154198,0.000796271436613649,0.000872375714834783,0.00785914875831506,0.000351865199652801,-0.0275061756106754
"2989",-0.00683670463082831,0.0011987901805961,0.00350883571233229,0.00604692073556601,0.000614097865898833,0.00208837207766965,-0.00174291348142264,0.00349538385361603,0.00826738808093386,0.00879950644204519
"2990",0.0104365506579378,0,0.0058888200471765,0.022288922775654,-0.000438171730708259,0.000694858007642685,-0.006235246969162,-0.00535898920978606,0.00113396721156644,-0.00186913334812067
"2991",0.00260063806455224,0.000239470960682997,0.000731778875828759,0.00195990237166344,0.00578728077879553,0.00307449677823635,0.0120466076966155,0.00377168080218038,0.00740616905304958,0.0062422403245177
"2992",-0.0169145298316905,-0.00766093339430129,-0.00438759533872923,-0.0134475129066624,0.00278988194334495,0.00148300859298067,0,-0.00214715223356643,0.000432407876689078,0
"2993",-0.0185061821643326,-0.017611560886834,-0.0183620576644139,-0.0215612706469214,0.00034770854844135,-0.000197359323472757,-0.010663356517672,-0.0134481825295959,0,-0.0303970519984572
"2994",0.00340754436098889,0.0135068501487652,0.0153385203672554,0.0184902351364764,-0.000347587689230378,-0.0001976331218001,0.00137869652735878,0.0111779279267255,0.00164262992379394,0.00831735623043794
"2995",-0.00667875533263729,-0.00799606190293978,-0.00368456684956497,-0.0116884552311891,0.00104339670673936,0.000592699979155453,-0.00337919184202973,0.00242645083001669,-0.000776834103427881,-0.0291878088056222
"2996",0.0161444144817968,0.0158768383911811,0.0134985447875449,0.0123300551167735,-0.0022582778549517,-0.000789903991447849,0.0035161634323162,0.00968258854723381,-0.00112289888026862,0.0045751006142738
"2997",0.00336436763483228,-0.00456834323410005,-0.000912262821317844,0.00695993319801302,0.00113169460834839,0.00098807627189279,0.00312860759849531,-0.000799111344238712,-0.00596681084371165,-0.00390365519694513
"2998",0.0230253903123594,0.0132848961015473,0.0131482500045177,0.0239447049662918,-0.00486912898272962,-0.0000987886678652794,0.00885733675337286,0.0130633070698596,0.00374075694843223,-0.00326592898342237
"2999",-0.00218504092596739,-0.00452921497374681,-0.00342458896192199,-0.0086788124346262,0.00393164994962758,0.00256621798545931,0.00136028415320499,-0.0115789864939716,0.00312013355313234,0.00655312555937493
"3000",0.00609528918470081,-0.00574710120540867,0.000904286720141423,-0.000972763366719254,0.00374263732560132,0.00196880366448937,0.00987882037674126,-0.0106497361690016,-0.00172798516896466,-0.00455729637804392
"3001",0.0132412048882988,0.0108381531861275,0.0135525519285171,0.0202044365046903,0.00710028185167544,0.0021858281236844,0.00464665713143386,0.00188363987293294,0.00752988568868029,0.0228908020595362
"3002",-0.0324022250133659,-0.0228734302016262,-0.0369048745983243,-0.0212359295611839,0.016741453976832,0.00461735363263216,-0.0154577208325442,-0.010475289518048,0.00609912357704245,0.000639377437478439
"3003",-0.00151720736628602,-0.0141429657793897,-0.00148103152358503,-0.00926389579246145,0.00314042518806912,0.00254249862806732,0.0250958604844962,0.0114007283219246,0.00017073086994368,-0.00830666140199077
"3004",-0.0232358946806729,-0.00964628591005889,-0.00741564119002847,-0.018700648237674,0.00186153728518912,0.00292620772685992,-0.0141101156867264,-0.00161038736490116,0.00810992836016666,0.0115979115668692
"3005",0.0018970335105839,-0.00774215340799289,-0.00765780097536473,-0.0105316944860415,0.00413822326822877,0.000583427626668964,-0.00562699360054342,-0.0083335230215712,-0.00347189443549467,-0.0159236109303792
"3006",0.00022712653820478,0.00352368123247637,-0.000752852132953397,0.00760268169370559,-0.000168188376004075,-0.00252701646316322,0.00073834524518479,0.00135546536608455,-0.00118965839564922,0.00582522978331501
"3007",0.00503544920692467,0.0175570181970115,0.0120549439894073,0.0163481605161597,-0.00445843508470634,-0.00272857833931395,-0.0164720064726714,0.00730909982304206,0.00212693549321985,-0.00321752554992527
"3008",-0.000338939189418852,-0.00172546592345701,-0.00297783832315668,-0.000247470171303332,-0.00236579039855045,0.000586466515349215,0.00599912032062933,-0.00322470083750004,-0.00220733506912862,0.0129115793058858
"3009",-0.0184647884779207,-0.0143209604945352,-0.0113869908236615,-0.0141089012930853,0.00347238486475909,0.00156241633169452,-0.00198761035809225,-0.00350502527664254,-0.00399898752658046,-0.0152963551974954
"3010",-0.0196184219935627,-0.009268400011339,-0.00793044969879053,-0.00928959883375968,0.00582383513277196,0.00292522723233235,-0.0369157095141026,-0.00730520591225381,0.00691957127831144,-0.01165045956663
"3011",-0.00109654056774466,0.000407424867303163,0.00278115775295884,0.00679082262430319,0.0059886608108719,0.00246459839576696,0.00897154777893494,0.00109020768362167,0.00237548988609082,-0.0209561733922374
"3012",-0.0149757111829021,-0.00687368299281554,-0.014728317287107,-0.016607005797675,0.0132109953109263,0.0034986163375017,-0.0109536442920404,-0.00490074874231783,-0.00609396519519312,0.00401346090748089
"3013",-0.016277862187858,-0.00410150083659278,-0.00524170709941196,0.0077942166101117,-0.00363107701029619,-0.0012591482379275,-0.0145928359958666,0.00136797965606217,0.0154134207613046,-0.0093271930529496
"3014",-0.020489685873923,-0.0123552580552218,-0.0308352539411487,-0.00696059900843082,-0.000165627469168039,0.00087291071927087,-0.0124287838750159,-0.0191256462506961,-0.00436092761423901,-0.00874238444107645
"3015",-0.0264228988331372,-0.0125097110629415,-0.0108740388359181,-0.00934579765737797,0.0049702726859866,0.00251881338757975,-0.0360157436771477,-0.00725830325740995,0.0109501009859325,-0.0110645613123692
"3016",0.0505248778800711,0.0250725569569386,0.0189332983323578,0.0199161525947584,-0.0107153560173747,-0.0047353287292472,0.0327779572276914,0.0187104439739849,-0.00299944183468026,0.0222376880571071
"3017",0.00767741592110105,-0.00411947972466886,0.0133866801414924,-0.00128464412761908,0.000166552084003957,0.00252458892906815,0.00161362543351662,-0.00367344112695389,0.00760484681247364,-0.00951735773123952
"3018",-0.00128998366696753,0.0085315489092963,0.00118281786591501,0.00951886617999276,0.00841383554089759,0.00542358772327978,0.00308830731739973,0.00226894572547165,0.00406401260678435,-0.00823610138714159
"3019",0.00875885261128362,0.00281964942742219,-0.00177229284042135,-0.00458705201958998,0.00379977825860922,0.00375696592401931,0.00307847411400264,0,0.00156948623111663,0.00276814258750346
"3020",0.00104026223999476,-0.0053680018445863,0.00690474164361232,0.00256015857204583,0.00526718337310172,0.00211128188674681,-0.0216172616417963,0,0.000659810309278308,0.00276057124542151
"3021",-0.0238628547339786,-0.00719602646791828,-0.00568182963944464,-0.0181307956022433,0.011379585727606,0.00794882387710483,0.00641006493786445,0,0.00906616650348369,0.00825877456338286
"3022",0.0334958058749315,0.0300284370333104,0.0338916293122373,0.0322495617634733,-0.0115752362811384,-0.00807595903101899,0.0107061270848989,0.0209394651155193,-0.00808623703340683,0.0136518996195234
"3023",0.00788467715740149,0.00150788931485679,0.00247750033611749,0.00226763981307765,-0.00294815101723378,-0.0027778666837236,0.0100565353115412,0.002771684274254,0.00345848973223828,0.00740742970686781
"3024",0.00939536705100941,0.00727722853754642,0.00475301027734654,0.0037707967194669,-0.00262836137211053,-0.00249749874279415,0.0181862492035834,0.00801551230077258,-0.00270804199320496,0.0100266691442319
"3025",0.00467345811406905,0.0122074025012044,0.0054871609271967,0.0177810629006114,-0.00156477137946753,0.000577882706220834,-0.00130371429636889,0.00740321191470494,0.00641816017788321,0.0198544006138881
"3026",0.00352752077840468,0.00147671458372667,0.00602184742025536,0.00713588151058797,-0.00643350659195419,-0.000480998455202108,0.0138382493142921,0.00653239187907984,-0.0058866978315214,-0.00259576096476599
"3027",0.000386350795822832,-0.00466945321738055,-0.0115974104349548,-0.00488650797614898,0.00390178673912889,0.00298459121367833,0.00347664529313452,0.00216335247084953,0.00172717334409644,-0.00325304643822777
"3028",-0.00610092828181341,-0.00419744636448527,-0.00359582565166827,-0.00834754282709316,-0.00372112642487576,-0.000575959164370698,-0.00320793748033721,-0.000270020909575508,0.00238089485104531,-0.00848568371229008
"3029",0.011460827151363,0.00223144510328099,0.0121557824182625,0.00693230276871293,-0.00365197667330619,-0.000960534594298901,0.00991239530395394,0,-0.00172003445720481,0.00790000123072776
"3030",0.00241969001510922,0.00024740644419774,0.00487890999653917,0.0122940762087345,0.000999551095163698,-0.000576914465651335,0.00624607563536084,0.00296912270604754,0.00319986880209711,0.00522536480298497
"3031",0.00758684614056726,0.00519414674543461,-0.00205420031271708,0.00437211730981124,0.000249515577364523,-0.00182766145633939,0.00532055230975281,0.00376752086229781,-0.00130854669113967,0.00064975053065397
"3032",0.0133099827814789,0.0125493212111805,0.0132860012400995,0.00483685024116043,-0.00524150641516774,-0.00318038162078582,0.0037802471238757,0.002948981002872,-0.00892641054027998,0.0103896539161537
"3033",-0.0135105182544555,-0.0133658319161766,-0.0179131270474027,-0.0173285249640331,0.00677473456881916,0.00348037948089175,-0.00288727352425766,-0.00534620117490536,0.0035531318018458,-0.00706942989049986
"3034",0.0020925217417016,0.00689661640216643,-0.00282072220544771,0.0102865739916451,-0.000415208280915347,-0.000481703444180082,0,0.00618128128818141,-0.00139973655166081,-0.00129445445557619
"3035",0.000531305007236638,0,0.0058457637791125,0.00969705048382363,0.00656540925892002,0.00318107468610074,0.00352498043416016,0.000801151041986747,-0.00156664744035828,0.00259226447945782
"3036",0.00846168654114399,0.0102739403546883,0.0108735858952851,0.0132052419545243,-0.0047887544299271,-0.00230596137246797,0.0116673499047704,0.0122765702015997,0.014617268630515,0.00517138674472584
"3037",-0.00760042607274891,-0.00460048564748361,-0.0072328962943502,-0.0104267199382028,-0.000995487672372897,0.00028896221655117,0.00905244721242515,0.0058000884892242,0.00349991857805709,-0.0135048870193266
"3038",-0.00132691343644464,0.00316227536958258,0.000934144450564833,0.00167646762614693,0.00506597587535951,0.00288837100616379,0.00798827303981064,0.0104848829323478,0.00559657713037076,0.00977835680421557
"3039",0.0158307837243057,0.010669204021897,0.0111981575203395,0.0217546832104978,-0.000743731611950849,0.00230419609790511,0.00792496624560934,0.00804146311416098,0.00572672191337187,0.00710137726681648
"3040",0.00878247408587041,-0.00143958868636518,0.0018456659164412,0.0084229280480268,0.00860009724445643,0.00459765001941315,0.0105238367162011,-0.00205872129710782,0.000481177312035008,-0.00512816137458549
"3041",0.000481544895179153,0.00120141606343682,-0.00405297697601126,-0.00788862035819982,-0.00603978673607264,-0.00535068522717896,-0.00682324101484577,-0.00128923940174619,-0.00200400801603207,0.00902057392904099
"3042",0.00703527440047091,0.00287989336238592,0.0022197076907633,0.00163709156076131,-0.0044642640790048,-0.00220934283412078,0.00674948622316118,0.00206563146751204,-0.00433735742971886,0.000638547936024469
"3043",0.00419195172570785,0.00909288585172496,0.0040605334044217,0.0137753317300862,0.00456725396196345,0.00173292288050475,0.00610576789189143,0.00154620368597524,0.00258147791692065,-0.00446711284627554
"3044",-0.00131826213942088,-0.00450547515457422,-0.00827205016349652,-0.0135881504500385,0.000495928652615163,0.000768522002423611,-0.00690165277294186,-0.0061744286865838,-0.00675890736046758,0.00128200777892928
"3045",-0.00953270829777231,-0.0131014726676126,-0.0139017652922642,-0.0100396690304838,0.00661009071382046,0.00326535824187624,0.0076683074271755,-0.00310638001972363,0.00243029808116813,-0.00960307277514072
"3046",0.00122154947100683,-0.00362057510128089,-0.00883458233863199,-0.00566046828613409,0.00426815971977224,0.0013401067250034,0.00023793296828778,-0.00103877404483266,0.00379829487309347,0.00129284668618146
"3047",0.000554400361612029,-0.00242244529859437,0.000948180270546439,-0.00332068151629605,-0.00392302591487459,-0.00152948400945219,0.0028529982629466,-0.00285938016550047,-0.00491104584905433,-0.00581019987504727
"3048",0.0128594644603943,0.0109275893619649,0.0176203592499558,0.00832933831836313,-0.00254361944644244,-0.00134044200921302,-0.00580840724902298,-0.00052153514183706,0.00210358417643342,0.00584415558710938
"3049",0.00324691994264126,0,0.00242037905314807,-0.00708039449859676,-0.00378424508579367,-0.0024923677726324,0.00465008171290227,-0.00756381843660692,-0.00395606326533127,0.00581019987504727
"3050",-0.00221820652335281,0.000240215423986001,-0.000742875014241973,0.00190159858436378,0.00569767432148938,0.00470914770297637,0.00320442329437021,-0.00289109012230748,0.00559289116658279,0.0025673722456947
"3051",0.0108972816071724,0.0158500838956881,0.012825249438412,-0.00142350430684635,0.0015602469813687,-0.000956602002169404,0.00615175284270308,0.00711649212989895,0.00596489611421736,0.0185659623806202
"3052",0.0017305445969249,0.00401900503876074,0.00165171899852168,0.00784029931851804,0.00254119858353441,0.00172346543482238,0.000235089074610118,0.0036641086404452,0.0152243105314669,0.00251418451559937
"3053",0.00201556017364268,0.00565092091284569,0.00109931764273763,0.00565770238089724,-0.00286197081349993,-0.000191231077810161,-0.0070530245182806,-0.00260774098544003,-0.00173633784695348,0.00313475350515446
"3054",-0.00355579249000515,-0.00468272525616531,-0.00146414729403155,-0.00210964469700015,-0.00893877602355042,-0.00296355820708427,0.000828598975888495,-0.000522682813473674,-0.0113061350891966,0.00312495753357278
"3055",0.00619975955963836,0.00305822941846268,0.00219936578929025,0.0110406920171999,0.00595776109464352,0.00297236698967085,0.00532292544629676,0.003138882531734,0.00359853649903541,0.00249225404025921
"3056",0.00136148781997947,0.00211065595336479,0.00566936428893228,0.0111523066558934,-0.00296130186817989,-0.00152956163408591,-0.007295006194322,0.00104310810725328,-0.00103583266932272,-0.014916033180699
"3057",-0.000715533647491662,0.00725487998612651,0.00345516123424439,-0.00344672008236058,0.00495006270042531,0.00296809809605825,-0.00272609020746806,0.00442825355766496,0.00167503385957479,0.0044163819462697
"3058",-0.00042978227264634,-0.00348523716416482,-0.00525553796897271,-0.00853120480077851,-0.0113289968492372,-0.0035322272017938,-0.00285232030016458,-0.00440873058078584,-0.00708711566989773,0.00502508265366841
"3059",-0.00186256746839164,0.000932682843835408,-0.00965560986849379,-0.0130233456549481,-0.00340432484005793,-0.00258660081749418,0.00297968533482273,-0.00468894898846839,-0.00561395451737989,-0.00250004222829769
"3060",0.00624394034079834,0.00628936518390777,0.00294324527018675,0.00117826576372226,-0.00924308883272917,-0.00328150055321552,-0.00213898283677616,0.00209386033736414,-0.0170175097510687,-0.0112781954887218
"3061",-0.00363738374525857,-0.00416666384170594,-0.00311810477133323,0.00141208924674929,0.00783744096534589,0.00308952205956436,0.00416811711115583,-0.0036563645537615,-0.002625525171288,0.00316865365604024
"3062",-0.00136022072075015,0.00209198799672161,0.000919974873967444,0.00987083239988085,0.00209052561874334,0.000577538203303751,0.00308344330461274,0.00550471807957464,0.00131624714241929,0.00505365229360066
"3063",-0.00605670504067868,-0.00185577339983056,-0.00588229506850624,-0.00558545378861086,0.00367147306685922,0.00278985795154796,-0.00484743019862988,-0.0059960879155726,-0.000903713433259012,-0.00565681936947671
"3064",-0.00836566692795004,-0.0146408062274235,-0.0118344498216857,-0.0184880658792506,0.00648475597074394,0.00335753788334436,-0.00178210391486533,-0.00131101082692786,-0.000822292567862037,-0.00252848771387459
"3065",-0.0019999008721745,0.000707534334004833,-0.00168407617001021,-0.00715315985792553,0.00421290442905464,0.00143431457318854,0.000952060135529953,0.00709020871740162,0.0109455516262769,-0.000633692099297978
"3066",0.0145013028935617,0.00848455691762418,0.0108716248781064,0.0187319863950874,-0.00296120151513068,-0.000763713511835462,0.0147444145113333,0.00547598081210521,-0.00488438635247102,0.00126825226655392
"3067",0.00377098158806644,-0.000934862395525538,0.00241058180313347,0.00518623734985946,0.00701251952143278,0.00277078441823808,0.00410130371936268,0.00233390535211297,0.00605370592365362,0.00633316485474422
"3068",0.0066192530936855,0.0109941900464547,0.0038844884588356,0.0011725691548039,-0.00188426435246736,-0.000381058479489216,0.00455121828632299,0.00569230206449967,0.00699294990259514,0.00629318041424543
"3069",-0.000639936342141878,0.00439611403626827,-0.0106872693329787,-0.00538764152939908,-0.00722319969311991,-0.00142993928073742,0.00151028534284858,0,-0.011547093396224,-0.00437765136383261
"3070",0.00494070517829126,0.0110573045343649,0.0115477480556092,0.0146020860903104,0.00661448352623983,0.00315011476033433,-0.00231988301259856,0.0051451598173502,0.0045747649840775,0
"3071",0.00362582492034558,0.00455692333696245,0.0027619573670068,0.0111419516501148,-0.000575084440599616,-0.00133218168086968,-0.00558068535572476,0.00295659729088626,0.000569244526557489,0.00502508265366841
"3072",0.00024793137724255,0.0036289541372112,0.000367189965442272,0.00045915017722975,-0.00221876639158258,-0.000666906086391306,-0.0029229856884021,0.00179464181546396,0.0027632964664881,0.00250010572949733
"3073",-0.00301001043000226,0.000225897925341556,0.000550667794275039,0.00160635934935582,0.010460126698475,0.00696036147364065,0.00334209845916966,0.00614111947671647,0.00648405754135339,0.00748116896669782
"3074",0.0112948472691143,-0.00271120278178338,0.00660432006854528,0.00137449167688031,0.00220106702624001,-0.000473584236158175,0.0169491307993352,-0.000762897674842389,-0.00402641327105813,-0.00495051590324702
"3075",-0.019246246361266,-0.0228816972679566,-0.0107527119723249,-0.0292840091311235,0.0155347933076915,0.0073892654146559,-0.00601852810973669,-0.0106897177419757,0.00234476875808531,-0.00870642553817436
"3076",-0.000752108252824457,-0.000463794871844669,0.000552696778389095,0.00235681846608626,0.00160180231175455,0.0025390104008769,0.000232854836291319,0.00643159858090558,0.00766312004788983,0.00376411527292286
"3077",0.00745413930269567,0.00417545981899137,0.0110477157604367,0.0030567062564455,-0.000719764522813082,-0.000844267138393917,0.00745066928228422,0.00409001782908147,-0.00496313648676172,0.0018750634218232
"3078",-0.00522916619774771,0.00207896435162214,-0.00346019522443164,-0.0107828360468262,0.00920231897126089,0.00291022959263132,-0.00208007370693852,0.00127290472138508,-0.00522929190918853,-0.00561453565263736
"3079",0.00379041441656991,-0.00437999608638262,0.000548252554077644,0.00663496911492722,0.00348846823213589,0.0000936793546735259,0.00868455389969736,0,-0.014152850559598,-0.00313672023395206
"3080",0.00630551275360136,0.00463070695147838,-0.000547952137918473,0.0103578243909765,-0.000947905132180571,-0.00159122873222839,-0.000803676679751786,-0.00127128649480368,0.000902378984374508,0.00062924131247688
"3081",0.0118592000181383,0.0124453530666637,0.0126096394603703,0.0165423550361008,-0.0142041132254818,-0.0068764252534087,-0.000344567135398988,0.00305498271585858,-0.00393412828564654,0.00943396226415083
"3082",0.000489787292154986,0.00318691784262537,-0.00685799902867379,-0.00320861007007989,0.00184936510411227,0.00170281287671492,0.00643606796756035,-0.00456851733230046,0.00370282237885977,0.00249225404025921
"3083",0.00157374016261258,0.008168816608223,0.00599674910269465,0.0068980515357171,-0.00866784897696571,-0.00311625259187565,-0.0010278159905287,0.00382452763573315,-0.00147565170989539,0.00124302907589291
"3084",0.0026534223614243,-0.00135057921637405,-0.000541914385633224,0.00616582842624647,0.00283366141205765,0.00104197860292721,-0.00148611331670034,-0.00482591820981704,0.00254513951038238,0.000620774470232011
"3085",0.00483997626081178,0.00157769275736674,0.000722869880482424,0.00771666818747341,0.00129149499467918,0.000473116914103455,0.00686886531383957,-0.00765703530851225,-0.00106459748534438,0.00310163159940502
"3086",0.000762531979169312,0.00180023385315753,-0.00234772302281283,0,-0.00354735753041324,-0.00160790070325467,-0.00591218663754556,0.00282940808552823,0.00434496628107151,0.00371063797274185
"3087",-0.00512486559353054,-0.00539090252099572,-0.00543093445029197,-0.00202699270261641,0.00315576534254425,0.0018000064167516,-0.004803954935791,-0.00641211868611491,0.00522406325648417,-0.00184842871977575
"3088",0.00341107909728788,0.00338763817986965,0.000182019060857685,0.00473938066816149,0.00241963423724578,0.00236401860224356,0.00907931430028319,0.00877660204586905,0.00308564347404561,0.00864193295515259
"3089",-0.000277664574861447,0.000224982741944935,-0.00309370471950265,-0.0107817512516121,-0.00587389220089629,-0.00226407843485621,-0.00102501624012641,-0.00332662089414981,-0.012790431577677,-0.00489591927758426
"3090",0.00676598617761814,0.006300759640264,0.00511136306296778,0.00726621544633055,-0.00712259334173693,-0.00463322404065702,0.00524467269320494,-0.000513401097571031,-0.000983968863894291,0.00307492641515528
"3091",-0.000654996847366807,0.000894352366552109,-0.000181622356089539,-0.00518490814387518,0.00252701660105781,0.00133015132797487,-0.0051038704585723,-0.00411000772234626,-0.00188790935093308,-0.0018393001365179
"3092",0.000655426149428262,0.000223394146288136,0.00399636158321415,0.00747795914197891,-0.00626111579765287,-0.00341541692359759,-0.021431881399321,0.000773749128404111,-0.00896378304216749,-0.00368550360883424
"3093",-0.00244703258744872,0.00402057038182768,0,0.00292392167073974,0.000409230861829091,0.000190290116286018,-0.00908654797833053,-0.00541231564587974,-0.00190858016913809,-0.00369913679082623
"3094",0.00196936989975316,-0.00200218852141876,0.00144745822365699,-0.000672839343960341,0.00523470612810573,0.00237954253865036,0.00681870185490929,0.00155480333384772,0.00074828733578558,0.00309401742611271
"3095",0.000861802994120531,0.000445815632396096,-0.00361335950592456,-0.00650810566508708,-0.0048007725946303,-0.00142442566008905,-0.00980844855739871,-0.00155238967320848,0,0.00493537152270385
"3096",0.00899172863573883,-0.000445616969384943,0.00562099279845163,0.00225886166017286,0.00212588605471198,0.00180645759517351,0.0119102167549585,0,-0.00207692941571169,0.00122758060901673
"3097",-0.00221929236036145,-0.0055729635612235,-0.012261077916811,-0.0135225775650958,0.00815858221651555,0.00379680094413803,0.00652617068074002,0.00207310973877184,0.00291373619096569,-0.00367860027303579
"3098",-0.000615862697940561,-0.00201742504099167,0.00219060832670159,-0.00137079443052202,-0.00145661095057992,-0.00122918695690311,-0.00196836475862672,-0.000775836727594847,0.000830073870423442,-0.00184621621650349
"3099",0.0046566900637075,0.00134768451222023,0.00910754605103947,0.00388931206463727,0.00340373065616273,0.00265050903106112,0.00754078296707394,0.00258794715121846,0.00663517458737672,-0.01171384965108
"3100",0.00156765389747227,0.00471061785409477,0.00397103910562713,0.00205101341812641,-0.00638067578524415,-0.00207703553236582,-0.00955689775942037,-0.00154878326768071,-0.00444921303989754,0.00062387250715612
"3101",0.000510475638938246,0.0046885319716794,-0.00359581890405136,-0.000909808197073536,0.00512124018208238,0.00198700756486425,0.0113928286150733,-0.00258515538187665,0.00306211200757911,0.00311710095042761
"3102",-0.00751643264619672,-0.00755556648605615,-0.0034284086344254,-0.00751191041504529,0.00412503911533157,-0.000454292826070124,-0.00068972805340306,-0.0028513223888863,-0.00660061897526276,-0.0031074148247241
"3103",-0.00215898676818504,-0.0042543677026603,0.000362201179833654,0.00229357346209658,-0.00476189955949846,-0.00283992203903527,0.000345156296592819,-0.0122172498247209,-0.00382059794317935,-0.0112220701642258
"3104",0.00978780839495097,0.00966957940285185,0.0128505988667482,0.0118994227538056,0.00283837058427916,0.00132935067590711,0.00793357827753538,0.0202630750850943,0.0059196263811967,0.000630495656581909
"3105",-0.00411523932822011,-0.00913146246094498,-0.0101858109552787,-0.0205789815397598,0.00274935961912059,0.00255940826351564,-0.00330818206537997,-0.00412696959926884,0.00132611684498762,0.00315068397557128
"3106",-0.016699708045074,-0.0188806817085043,-0.0182343464264934,-0.0196259965445982,0.00766127623377022,0.00340425755513052,-0.0181983824915457,-0.00207192020842906,0.00331099252232425,-0.0125628342747678
"3107",-0.00138928336036537,0.00504005648486672,-0.00606842767564142,-0.001413013881988,-0.00432177626649233,-0.00188483772423187,-0.000116514275515622,-0.0028551098763212,-0.00247500208295515,0.00127222146063866
"3108",-0.00302566152528005,-0.00569860798348765,-0.00647545365394009,-0.0158019300682993,0.00409942996785229,0.00264401626675626,0.00233180334067051,-0.00025996531526129,0.00239842023328363,-0.00508254897919436
"3109",0.00502338108377165,0.00664836611589159,0.00689010264621115,0.00599077019595717,-0.00136081018851486,-0.000659321089255038,0.0105850217890313,0.00702924211873102,0.00189771456842536,0.00191564380807363
"3110",-0.0251303345622579,-0.0214074254542168,-0.0225632686190562,-0.0333490524573676,0.00785572135622803,0.00499447374993189,-0.00115109035558703,-0.00646319193435452,0.010211628098493,-0.00509874586703907
"3111",0.00904387394539441,0.00791243486394588,0.0140018156744555,0.0140462764762501,-0.00294279077675064,-0.000937867160224481,0.00414855830929617,0.00468371328109929,-0.00171190187840398,0.0134529142144599
"3112",0.0058573866649001,0.00600318851007975,0.00149275795174897,0.00194411309996045,0.00614223883006138,0.00319094417033083,0.00654106545866395,0.000518153783467978,-0.000571615225964495,0.00884951432741188
"3113",0.00926127312513891,0.00895109595364163,0.00409919573086692,-0.00485082703871986,-0.00332988812338852,-0.00196441804744851,0.00592863835584434,0.0056947718951228,-0.00719010545951559,0.00563909774436078
"3114",-0.00646525114483332,-0.00636936764217122,-0.00371125345357015,-0.0180355019530282,0.00222717091083213,0.000468547996425261,-0.00283344478500436,-0.00669220069517351,-0.00707760666484059,-0.00934579439252337
"3115",-0.00661191722912391,-0.00663923390975363,-0.00540131253522147,-0.00421955714561073,-0.00206344094635125,-0.0016865283372659,-0.0147760555853503,0.00492346180819681,-0.0000829092402335752,0.00440255832365777
"3116",0.00901557495446603,0.00691405557179747,0.00692873354950518,0.0127119247539218,-0.00159074753544364,-0.00112606953502148,0.00842179894226458,0.00361013869264415,-0.00232093834815106,0.000626152843005601
"3117",-0.00307150480673934,-0.00389104424870801,-0.00818291426398265,-0.00492256309267958,0.0057355392466667,0.003006365290946,0.00354641020367286,-0.00693724853411204,-0.000997033890021259,-0.0143929485468923
"3118",-0.0122185484719306,-0.0101101757938219,-0.00750052485030617,-0.0128617526345564,0.011247629550396,0.00608924636141617,0.00136803818378439,-0.000776122523459155,0.00773453106677535,-0.0209523796007606
"3119",0.0022683797064289,0.0106776714490011,0.015492122526958,0.001002362101163,0.000861794071915778,-0.000279367792606511,0.00330130715824217,0.00828576522543956,0.00107291410535471,0.0136186761454711
"3120",-0.00930052004639614,-0.0105648633096769,-0.00837202713387675,0.00350437862068387,0.00719969916908214,0.00437752216799381,-0.0105525030827032,-0.0118130951388754,-0.00387469899732817,0.00831731624288978
"3121",-0.00671067457374919,-0.00928520618013995,-0.00469043291453963,0.00648541547723025,0.00303038934892941,-0.000371005279576897,-0.0119265291729143,-0.000779580448413975,0.000331051885607003,-0.00380710643535986
"3122",0.00273125094500881,0.00585759427031318,0.00452403295378545,0.00545229685341853,0.00859846488757987,0.00361784096952267,0.00406213043268999,-0.00182054683686317,0.00678413981672543,-0.0101910607913405
"3123",-0.0134753266845519,-0.00931757714778059,-0.0106961328288799,0.00345082387176099,0.0125195146574724,0.00665488641723377,0.00416140909514806,0.000260556628771891,0.013476867228583,-0.0263835464521808
"3124",-0.00254311873671986,0.00705398812971425,0.00588000021162749,0.00908871107116971,0.00668885123915164,0.00481150224173832,0.00391387794076925,0.00859615809224268,0.0144328141663372,-0.0033047148998443
"3125",0.0217068443455004,0.0121408352915391,0.0115028750200419,0.00219070908637686,-0.0114013934221635,-0.00366231288277741,-0.00321064809293237,0.00413206723473247,0.000319726638000839,0.00596816962723756
"3126",0.00866215128486014,0,0.00055929125280052,-0.00801550230660464,-0.00565183047261419,0,0.0209364622585657,-0.00411506351561075,0.00255692365070836,-0.0204350464341544
"3127",0.0065026396519714,0.00553649835246439,0.00111803395091314,0.000489806251149361,0.00322579643575205,-0.000183683343144336,0.00146468180765158,0.00335708808101054,0.00326768149145074,0.0174966572558402
"3128",0.0100069599807269,0.0126175685106944,0.012097505436762,0.00783154333565017,0.00865178022560609,0.00395224585028897,0.00303778915045294,0.00566310063342224,0.00564028453225962,0.00330683328664261
"3129",0.00458894472269056,0.00203893003913147,0.00459727992867132,0.010442014435319,-0.00941232541406389,-0.00494382059804255,-0.00302858893584246,0.000255955010062703,-0.00995334576043438,-0.00263676074053543
"3130",-0.000242230813356836,0.005200059626562,0.00329487817278151,0.0112953164582721,0.000612999512164647,0,0.00168760561463155,0.00511761863525617,-0.00119685628027033,0.00660936264706513
"3131",-0.00176517678752663,-0.00584791056377054,-0.011129403343153,-0.0106938829005175,0.000765760374777491,0.00257614321502153,0.00325736974814528,-0.00865583179715668,0.00519253874420822,-0.0137885081622434
"3132",0.00412613724282251,0.000905039914101513,-0.00110694921685317,-0.0016815285357209,0.003443480732221,0.00247759801198644,0.00369463787894331,0.00308165702068619,0.0061193355142759,0.0126497765772546
"3133",-0.0011049433468322,-0.00791147755600186,-0.00258586419461238,-0.0110683331395599,0.00251669137438126,0.000732421868165023,0.00167311078564669,-0.00409632910581226,-0.000315955771184151,0.00394477291203388
"3134",0.000380411623847055,-0.00046768047406498,0.00293378139210709,0.00394713031967453,0.00174956794631043,-0.000182992436909557,0.0107165053802742,0.000514175993955979,-0.000632071754615549,-0.00458419598484128
"3135",0.0104709756119306,0.0142722282152554,0.00596241036073608,0.0241759138802855,0.00501186171612478,0.00192140383639261,-0.00177621054223764,0.00668047936755345,0.00506008843152861,0.0118421049993025
"3136",0.00225708951169157,0.00438300083078125,0.00889056831585666,0.00834522424872297,0.0014355253610383,0.00273945378992946,0.00622835399453603,0.00280754347008538,0.00605723711318662,-0.00195051907153276
"3137",0.00955431653183436,0.0101056076693329,0.00973011257376255,0.0146606648234773,0.0026406042729803,0.00163921151927138,0.00442136412488581,0.00763562648919791,0.0251779030821637,0.0201954158937032
"3138",-0.00145362363823298,-0.0015916254368471,-0.00981816247769951,-0.00326261165311603,-0.0109866465762964,-0.00409121566670723,-0.0126554288032473,-0.00303106101932626,0.00663561126812895,0.00255425662399422
"3139",-0.0012243298597332,0.00159416274682544,0,-0.00140286993750149,0.00745644897193576,0.00346883998886427,-0.00624162537851825,-0.000282025293394716,0.0148507808713678,0.00445857696222429
"3140",-0.00980814852358014,-0.00568438318078257,-0.00440688289700653,-0.0103020692628075,0.00309652782659797,0.0015466533652968,-0.0127860999150258,0.00102514813054744,0.00194113032789112,0.00317059845271306
"3141",-0.000997215153538344,0,-0.00147546315902958,0.00946294861205321,-0.00639966839335071,-0.00408764787803917,-0.0188592933046174,-0.00512040648066303,-0.00916539513782555,0.0050568469803165
"3142",0.0035459176287056,0.000228734864551106,0.00406354751927873,0.00703086105453377,0.00704718348979649,0.00300996335388337,0.0115794042847437,-0.00257332309398028,-0.000977701729880986,0
"3143",0.00514581202430509,0.00754454393708381,0.00404708316520042,-0.00139643591952299,-0.000677253542837208,0.00045470753285648,-0.000572290444978085,-0.000257870718607278,0.00271003470972686,-0.0106917812989837
"3144",0.0090784728658817,0.00294989534628587,0.0142908891068925,0.011885310246645,-0.00233847499578899,-0.00125652579388325,0.00343605432469452,0.00335475316468092,-0.0193693848206319,-0.000635706350688436
"3145",0.00260435036327289,0.00316733720484841,0.00307086362908437,-0.00253331998948569,0.00771282272959617,0.00355559741667544,0.015637456939694,0.00488692362148435,0.0213597389894249,-0.0165393960464058
"3146",0.00799507778371078,0.00721695710836112,0.0028812379801475,-0.00184719516399534,0.00712914493258254,0.00190762127815702,0.0132614811229927,0.0133095578577602,0.00164905924146463,0.00970239117406657
"3147",-0.00113783165910819,-0.010747834525742,-0.00430947707668383,-0.00693959310311443,-0.0132631112083185,-0.00634697818625629,-0.004547531614429,0.00176783738934194,-0.0111502353083054,0.00192190997549258
"3148",-0.00549480311393369,-0.0045269708629494,-0.00577101041243011,-0.00605644626971125,0.00135936067421505,-0.00100363355873212,0.00323116687433966,-0.00352999281323829,-0.00643261697012709,-0.00127885885720846
"3149",0.00124649446826508,-0.00409275774393536,-0.00888801687440532,-0.00304659089620518,-0.000377135940662132,-0.000639262613443048,0.00488678355061767,-0.00328939031474451,0.00350374761616434,0.00320104594039505
"3150",0.00477809029937948,0.00365302477068252,0.00603955338781104,0.00846260832455958,-0.00550673960866466,0.000548340377880541,0.00530499045764921,0.0020310933994796,0.0157874914611007,0.0216975534556096
"3151",0.00234409021264281,-0.00159246536598789,0.00181915591477266,-0.00186475333630609,-0.0133507679387136,-0.00493287938641163,-0.0112137252112869,-0.000253540108381523,-0.00844358501914999,0.000624588412292182
"3152",0.00447705713967594,-0.000455616303364104,0.000363144589517805,0.000700555939275427,0.00115360412773713,0.00110151336355235,-0.00177903210380892,0.000760420992281352,0.00625472508488456,0.00249679418045523
"3153",0.000332418777221122,0.0018236211603242,0.000726044041240881,0.00373388247276063,0.0057592487448086,0.00210912870408109,0,-0.00202597789148029,0,-0.0105851998891362
"3154",-0.00322499606810767,-0.00341303655211644,-0.00743690830286692,-0.00139494641650717,-0.00297766275667954,-0.00219619464893517,-0.00233906719700205,-0.00304484167050523,-0.00846255529440998,-0.0106985729502709
"3155",-0.0068051869214466,-0.00205483515877547,-0.00091377086411315,-0.003026729432824,0.0107980240994714,0.00467726963638349,-0.00401923570742957,0,0.0164653179667065,-0.00890587338578497
"3156",0.00366107431359741,0.00503325739078275,-0.00256083506122196,0.00607200460815682,0.0000755632643583137,0.00246449931272386,0.000224399849312107,0.00432672091898789,0.014117951937614,-0.00706035519196246
"3157",-0.00555503537890945,-0.00614619328257104,0.00256740977418835,-0.00510679359716049,-0.00234833499893949,-0.00182094381459386,-0.0146812153088112,-0.00405470077845793,-0.0147273963870866,0.00581777724944499
"3158",0.00245640622424648,0.00206142420430977,0.00146331832925517,0.00023323678051268,0.00189847298340018,0.000455920207446558,-0.00181990606808224,-0.00559787626312769,-0.000148761804500963,-0.00321338909511093
"3159",0.00715015751186998,0.00640001766614517,0.00803652812536138,0.0011663193372855,-0.00545713896425115,-0.00164127001628267,0.0101413066867251,0.000511490024671657,-0.0056526219186156,0.0064474309978213
"3160",0.00469952945760443,-0.000681459647587479,0.00126827028768117,0.00163097359156916,0.0043435889418808,0.00146137427105919,0.00281997767400854,0.0015347317601031,0.00508634146029863,-0.00448428304224902
"3161",-0.00477707431016672,-0.0104544594301914,-0.0106767175337291,-0.00883927930291684,-0.00478043703345488,-0.00173284902498461,-0.00461181027070623,-0.00561803018370721,-0.00707000844943095,-0.00386106898946703
"3162",0.00669988146333877,0.00528254855108234,0.00256081640453854,0.0021121462682987,0.00236397486518181,-0.000182718364506562,0.0033902469088094,0.000513584552739532,0.00164893571651836,0.00129201154218861
"3163",-0.00182110959728077,0.00182771756658728,-0.00127713768712923,-0.00187348751843941,0.000304178818301137,0.000913842473360571,0.0029283027718443,-0.00359333156116071,0.00665968277955487,0.00387103320698201
"3164",-0.00245462120968398,-0.015051352390594,-0.00639387290072335,-0.00774287977732702,0.00243328858763503,0.000456327545628188,0.00718691055855047,-0.00644004998621805,0.00334495654013933,0.00578399589622292
"3165",-0.0109403776746063,-0.00648290576207167,-0.000735463264501579,-0.0122960344124852,0.00804039270861079,0.00255520843546231,-0.00334487573089848,-0.0111484238000432,-0.0131129726807816,-0.00638968965774234
"3166",-0.00870800016427153,-0.00419483768845952,-0.000183912001185282,-0.0196313867266756,0.0198603732473872,0.0113421982404234,-0.00100674783869958,-0.000524444055387652,0.0240221967708476,-0.0276527736668752
"3167",-0.00752941826821574,-0.0100633458720004,-0.00515275443678287,-0.00976798164921744,0.00924154126164001,0.00207368315034029,0.00447911740170515,0.00996838953012724,-0.0038120737830929,0.00132277363287803
"3168",-0.0300731777673868,-0.021749254506905,-0.0247872378782149,-0.0369913244791921,0.0172882741925715,0.00863694043017027,-0.0179487152137093,-0.0199999597990181,0.0139818530722045,-0.00858656973011873
"3169",0.0140229300208405,0.00410818979354621,0.0127085534066838,0.014340662391978,0.0079930587614867,0.00160568607146439,0.0105574679899101,0.00477087770665485,0.00812839144276589,-0.00532973477973142
"3170",0.0005907154823519,0.00505407984886452,0.00693013689789956,0.00454423359460376,0.000357232451593914,0,0.0104469970634213,0.00501184788790998,0.0151896907295461,-0.0127260991363837
"3171",0.019620099910866,0.010775905038946,0.00706850382829693,0.0123146891470816,0.00214240363185492,0.0000891120370902776,0.0167872059234333,0.00524922129272531,0.00503468997206946,0.00542736221015194
"3172",-0.00681161394504937,-0.00497505386851071,-0.0105282608007198,-0.0101788369260873,-0.00199529278000943,-0.00151380171349624,-0.000109399893315598,-0.00365525316394311,-0.0033161716874669,0.00877197552943043
"3173",-0.0121731653589806,-0.00785720079742036,-0.00952025053605543,-0.0120391231694671,0.0208498447190082,0.00633181478133982,-0.00382710664860209,-0.00445496034052772,0.00969849956457947,-0.00735781389097367
"3174",0.0155515948776324,0.00863928413446957,0.0113079175972337,0.0126936314675397,-0.00342755773271697,-0.00354481214408731,0.00109750008162357,0.0023691566436157,-0.00595951742412126,0.0235847893992234
"3175",-0.0295676261918925,-0.027123487103055,-0.0242266188168268,-0.0288291888139194,0.0225295124813343,0.00667032198168194,-0.0162279148995914,-0.0168067648948103,0.00684159265652129,-0.0151414293457932
"3176",0.0026417847073803,-0.000244422185778359,0.00954929648799174,0.00671130670751197,0.0111195343010746,0.0063608503362993,0.0110343282962551,0.00988250618086628,0.00665497022767081,-0.00802138964796029
"3177",0.0147550644352292,0.0119862214594069,0.0104047975132557,0.0138461946539619,-0.00801034464464512,-0.00263371829354297,0.00870902759997527,0.0134885086323775,-0.00640221307729039,-0.000673900029193431
"3178",0.0120476617952245,0.00773497199107265,-0.000187148797616721,0.00404642952205281,-0.0143024929005783,-0.00475305596134912,0.00754104200532324,0.00287050372352216,-0.0116963020849999,0.00472013878150723
"3179",-0.0076624856960561,-0.00575669496050846,-0.00205995803644166,0.00201516446386063,0.0103446000814065,0.00442205363528503,-0.0074846003199176,0.00286220121468705,0.00779537943593356,0.00268454096763349
"3180",0.00813533402518729,0.0118213940019076,0.00337777592674482,0.00955247734455278,-0.00666547374479087,-0.00264146880703919,0.00371584496729249,0.00337326291847306,-0.00316441866147987,0.00334674288307091
"3181",-0.000307756373121859,-0.00214586815164985,-0.00149623509115548,-0.0129482159866834,-0.00664080878494444,-0.00220726164318208,0.00555317250375942,-0.0036203931307186,-0.00253951052975143,-0.00466975715446305
"3182",-0.0256874733296693,-0.0126642032181168,-0.0112380247244338,-0.0148838701789102,0.0164346951315082,0.00672469110343998,-0.0137520167131248,-0.00207631314454215,0.0195898452442651,-0.00737260842225429
"3183",0.0110585038226301,0.00701837524838678,0.0145860398170012,0.0053777220900284,-0.00404221634512969,-0.000966877905066776,0.00735611464912456,0.00520152547181318,0.000138752863130476,-0.000675265120282376
"3184",-0.00392356925283832,0.000480703997335352,-0.00317399052335154,0.00178302051713874,0.015408701020307,0.00431076209650905,-0.00381469484005525,-0.00051732366381041,0.0095707398630871,0.00675673356420781
"3185",0.00704150277402493,-0.0007207462683535,-0.000374571531394419,0.00279673826879767,0.00128741435094337,0.000350324579709627,0.0022976087844262,0.00232981963944945,-0.00281653486490541,0.00872487747592454
"3186",0.0127729420240308,0.0100961822895875,0.00712008009091547,0.0111563263831447,-0.003788889442081,-0.00192643956169825,0.00796859754885482,0.0005163597825939,-0.00716456993208681,0.00266132126566654
"3187",-0.000444342179129475,0.00356970227742948,0.00316277075432159,0.00777322307773654,0.000271482786295296,0.00026322968239012,0.00129947679334141,0.00438829118585726,-0.00256727041934735,-0.0159256794434508
"3188",-0.00584719951049739,-0.00308268435181769,0.000556419720665113,-0.00622044105756414,0.00129263127433354,0.00219653492034122,0.00973401248103589,-0.00565423990284786,0.0139130434782608,-0.0053944247471307
"3189",0.0113505298840004,0.0164129728960816,0.00556070588025337,0.0167751533805764,0.00149430323589361,0.00157777788842006,0.00781905048105913,0.0129234080646554,0.00624359519725548,0.0237287654582146
"3190",0.0128552195358529,0.00514850222278529,0.00718898529457035,0.0113272489242768,-0.0181102881253071,-0.00805247305642776,-0.00627049508931365,0,-0.0240011243965328,-0.00132452568052432
"3191",0.000772418139330933,0.00209550132070402,0.00347725639413632,0.00438279088479532,0.00711512632284217,0.000617683272586156,0.00192514372063224,-0.000765547010674106,-0.00852313125976756,0.00265256475118081
"3192",0.000503292242964193,0.000464637945744695,0.00656575421803041,0.00315156688527019,-0.0177652337927561,-0.00617289454687675,-0.00651155260277825,-0.00229817471751481,-0.00373449131531134,0.00925928103607609
"3193",-0.000234857334677541,0.00139343214340948,0.00289906192241984,0.000724860374757164,-0.0175278259971099,-0.00727582347608957,-0.0106371433588983,-0.00307145166505018,-0.00855793202176902,0.00131050490558815
"3194",0.00711099286826733,0.00533390755234597,0.00885276325103845,0.00700318994819615,-0.00177699068818027,-0.000983318155923008,0.000977416042232226,-0.000256839854801516,0.00606367557744147,-0.00719890871020412
"3195",0.00346393376887,0.0059977572031471,0.00662607451165154,0.00719430982550961,-0.00655082212276048,-0.00223668620336426,0.00488231944819328,-0.00154078204874075,0.00205635681809802,-0.00395517459858208
"3196",-0.000663839906607233,0.00275164671388417,0.0117415991357641,0.00571423441982466,-0.021358932341752,-0.00914630189813337,-0.011660552635918,0.00823057378409597,-0.00827917451207039,0
"3197",-0.00308891358734265,-0.0107477653838878,-0.00527510125448916,-0.00781251235012204,0.0127436663410869,0.00434398527554958,0.0102687856011461,-0.00433676714081166,0.0083482914740618,0.0443414722905136
"3198",0.00253209353421213,0.00485437064741379,0.00371221055656834,0,0.00542354314497029,0.00261286303553265,0.0109210538656281,0.00614908562765315,0.00198131181807826,-0.0190114068441065
"3199",0.000598089146846226,-0.00092015394556022,-0.00211344595177188,-0.00405625149827993,0.00424369069249342,0.000359581097637118,-0.00352948185928381,0.00050926866148715,-0.00628530340599009,-0.00645992644230764
"3200",-0.0000664286097289413,0.00345390194241224,0.00741266422455689,-0.00407284551923504,0.00300807052750929,0.000449271528025319,0.00483026737438763,0.00610839464331847,0.00405082774247889,0.00520164843502324
"3201",-0.00472476134058997,-0.00206520813904432,-0.00227752553837912,0.000962194927357496,0.0132107916390476,0.00574706216257148,-0.000427448943598474,-0.000758962528595308,0.0118204842286274,0.0012935513870731
"3202",-0.000234757365234373,-0.00252931227273578,-0.00105350591466302,0.00096139344055679,-0.000211739222357954,0.00142856007074221,0.00149623870242244,0.00104781563549827,0.00559638346826974,0.00258408871869475
"3203",-0.00784666805641099,-0.00576300490134163,0.00140621570865607,-0.0105642579646796,0.012054412452071,0.00499281412986585,-0.00124659716662079,-0.00357407606328586,0.00528692173913048,-0.0115980023440451
"3204",0.00591474757755983,-0.00486912019834607,0.0040371437636213,-0.000728050012543724,-0.0146269890362218,-0.00656488227773222,0.000753145456512394,0.00358689590207084,-0.0185453815841596,-0.00586701408252943
"3205",-0.00208322105157543,0.00535885784137768,0.00174821664641178,-0.000242851836431579,0.00643233036363355,0.00214328170783862,0.00817211658941108,0.00638239051935185,-0.000282091232008841,0
"3206",-0.00538718764883572,0.00046345347114185,-0.0143105511369014,-0.0128734504453801,0.00245817360411205,0.00142568712180746,-0.00607933974833275,-0.00329770968614373,-0.00514842397939885,-0.0039344926789654
"3207",0.00463772560448916,0.00231652440461971,0.00460342230108379,0.00565948171602315,0.00245235967632995,0.000800960159485609,0.00375576395868316,0.00585379047943335,-0.0155253298670827,-0.00987485104181107
"3208",-0.0118947719856339,-0.0108620939960015,-0.00440601884770475,-0.0070956195021642,0.00301052645248268,0.00276942540858927,-0.0105837595255662,-0.00657903542414928,0.00547281650006548,-0.000664871068921102
"3209",-0.0176645964736546,-0.0261681781457669,-0.0123916664018512,-0.00763933875937273,0.0024428108996748,0.00346321663659044,-0.00388967270908658,-0.0056035309257545,0.0116736370524373,-0.0086494124123877
"3210",0.00819269446573423,0.00695785369340229,0.00501881470485643,0.0129128471844888,0.00912208616087051,0.00522117469803707,0.00976232136881827,0.00768443375981476,0.0045306457783747,-0.00134230457842133
"3211",0.0135321104459509,0.00905391607056449,0.011592664532686,0.00441297713061184,0.00738329021642037,0.0019368668349804,0.00537123298268538,0.0119471679895657,0,0.00806451612903225
"3212",-0.0043147139714127,0.000236212400573477,-0.00634690100736257,-0.00829880793602045,-0.00828806679508054,-0.00333886337510625,-0.00277804993549857,-0.00326540326940861,-0.00852707576576783,-0.0013333559115386
"3213",-0.0155246751496994,-0.0110953673366143,-0.00585525572016421,-0.00713753288462238,0.00269367352773098,0.00211580897380292,-0.00514310741410884,-0.00302425675985984,0.00874259707523506,-0.000667466324014487
"3214",0.0094964130167714,0.00811644481315277,0.00874526807231724,0.00768466092632125,-0.00564866124306862,-0.00255122246555317,0.00323106538221962,0.00505540397983828,0.000916044263191251,0.00267198788324197
"3215",0.00676344987545741,0.00899836749161498,-0.00123849821255106,0.0103320294834623,-0.0148942595517173,-0.00626224294132616,0.00193238666458995,0.00100617687383031,-0.00872935567625432,0.00666220231940717
"3216",0.0103668393511498,0.0211217889898547,0.0124003760611322,0.01607017488041,-0.0123767919954828,-0.00683409122429313,-0.000750094584719863,0.0100502516710979,-0.00553937228235746,0.0119126403683329
"3217",-0.00111367547379704,-0.00436688290357135,-0.00437442763282747,-0.00431349724283137,0.007262793644917,0.0027704681963201,0.000214484686451133,-0.00124372325531197,0.00399912164535543,-0.0045781334059144
"3218",0.00990034011688823,0.0129271853765356,0.0149385192136162,0.00890485967803967,-0.0120880828499514,-0.00481245552261722,0.000536057986276983,0.00697381249166518,-0.00697058843361797,-0.0026280985247561
"3219",-0.00160607469256657,0.000911556280349668,-0.00207801790962947,0.00286270492471163,0.00121631125706201,0.00197003217313263,0.000749928622351348,0.00692559650910662,0.00573026999691795,0.00131747834751383
"3220",0.00294908450918552,0.0047814222548892,-0.00260280301127591,0.00380592213810171,-0.00243000122141801,-0.000357470249887304,0.0055674028381405,0.00147372229113985,0.00142437856493483,0.00394743517647012
"3221",-0.00437720011691334,0.00067975378017926,-0.00191368663907421,-0.00521338367883073,0,0.000894022362129432,0.00798562690726357,-0.000245218646040102,-0.00106673777777744,-0.000655352323614466
"3222",0.00677914065107199,0.00407607526089504,0.00714655345035253,0.00905204312412899,-0.00752251248158942,-0.00366230984429183,0.00728848043453589,0.00588824938058319,-0.00477014072767334,-0.00131149755965509
"3223",-0.00326673437517733,-0.00405952831794731,0.00121156110391407,0.000708090725924926,0.00584690918776865,0.00233104734375944,-0.00325077555440434,-0.000731796062110823,0.00293299964611915,0.00131321984427624
"3224",0.00290967327787284,0.00634057433789104,0.00414864023169015,0.000236089415121876,0.00100498841306962,0.00035768552844484,0.00136760752509302,0.000244021558685859,0.00235379462953911,0.0124589936319914
"3225",0.00163401713169131,0.00360041597346172,0.000516406788504398,0,-0.00200751462174353,-0.000178842198316431,-0.00126086141989701,-0.00390432776182037,0.00711591835989411,0.00518143477574506
"3226",0.00409494797956977,-0.000672659009318899,-0.000516140250175323,0.00707536547001553,-0.00488514764067438,-0.00214620047071112,-0.0102041040233279,-0.00367473984778377,0.00233167527966982,0.00579890297429775
"3227",0.00563652360631428,0.00426284313198222,0.00292640463181981,0.00585478983729781,-0.00909631884842976,-0.00376404695113319,-0.00542024053404566,0.00122945804967856,-0.00860004223459732,-0.00384362468784738
"3228",-0.00029672048613949,-0.00134034980923758,0.00429120667391336,-0.00512227525287223,0.000656170916757404,0.000899425938652554,0.00341960070171687,-0.00122794833870898,-0.00277303045202659,-0.00192926024006812
"3229",0.00306727275434437,0.0062639080447191,0.00273450977307665,0.00444659245918455,0.014633897063163,0.00485361137971907,0.00553768000060795,0.00442591972660566,0.00549022459893056,-0.00644334190948614
"3230",-0.00266339675028504,-0.00333479085711863,0.000170491856401833,-0.00792166999326216,0.0134901709137882,0.00635047151222268,-0.00169445811134017,0.00342719556542281,0.00999850347472697,-0.0058365754909161
"3231",0.00926402061024922,0.00736112849222592,0.00988413049270154,0.0150304521321705,-0.00307811103462341,-0.00188700163723865,-0.000742617250360733,0.00390337517356243,0.000912764209712646,0.0182648168799422
"3232",0.00401766465361564,0.00465022485662603,0.00674986582677617,0.00994921014300654,-0.0131614976063804,-0.00508340692650444,-0.00775026920805477,-0.00121501033573157,-0.0028760101413583,0.00640612793002915
"3233",-0.00110618262090545,-0.00264497163380673,0.00134099392511189,0.00572736545801722,-0.0112465961184111,-0.00537824129283726,-0.0162637092561762,-0.0036496783116462,-0.0161800077177632,0.00254619201042838
"3234",0.0002279674656811,0.00132599303085668,-0.00217609868987279,-0.00318922261411747,0.00605147470834866,0.00288389901433583,0.00293664904698199,-0.00293027734405138,0.00429024650882015,-0.0107936716004128
"3235",0.00351686591026135,-0.000220781156841099,0.00587143972091853,0.00731272957699525,-0.018118447274863,-0.00799776940744235,-0.00954326705189812,-0.00269424542875596,-0.0155214884055853,-0.000641891971205011
"3236",0.00246616760580531,0.000220829911924625,-0.000500301395400471,-0.00907447648335635,-0.00420711478541158,-0.00135886587669365,-0.00186143691329299,-0.00982318329241527,-0.00636439556333568,0.00256908653475652
"3237",-0.00190982174417442,-0.00154492829065811,-0.00250292930292262,-0.00709705256125137,0.000666896336154243,0.00108857009018148,0.00230368029607098,-0.00471229439952836,-0.00240192883326229,-0.00640612793002915
"3238",0.0021078792914957,0.00110527597681265,0.00217465976164366,-0.00645603786195537,0.00459283215040185,0.000453029563051377,-0.00700455514768583,-0.00523302784300372,0.00269951120238598,0.000644788954934805
"3239",0.000323661301079747,-0.00198723273734736,-0.00350527077697904,-0.00765840137370843,0.00648881541681079,0.00271716631221852,0.00815594007556619,-0.00551099646610509,0.00400205943399845,0.00193298947981591
"3240",0.0014557539726352,-0.000221295908388486,-0.00435513064435189,0.000701538957995185,0.0103296420802659,0.00505816254456137,0.00798083798708538,0.00428214854773112,0.00420352237146027,-0.00321552085191401
"3241",0.00723653057534279,0.00464713768017555,0.00588836977002538,0.00794583319048781,-0.00108790821749727,-0.000808804268603636,0.00531456650636941,0.00777521560686112,-0.00252591660689849,0.00516131205968251
"3242",0.000737608500204434,0.00132152212088221,0.000836217791993388,-0.0016230323781169,0.00181486311704804,0.00170890833484094,0.00517853037961014,0.00746640862929393,0.00296641327859848,-0.0102695541958202
"3243",-0.000288522777752376,-0.00131977800505378,-0.0031751567248175,0.00209016874202406,0.00833285576578313,0.00188566672307156,0.00128798500652483,0.00370557784018444,0.000505028152684606,-0.00907920528324691
"3244",-0.00371870674387498,-0.00594718625466162,-0.00301751125017768,-0.00440338259509332,0.0103477794883589,0.00367463098300713,-0.000214415711430438,-0.000738352491468697,0.000504672283442753,0.0130890276901821
"3245",-0.00160899083110411,-0.00177270679627861,0.00100879564011769,-0.00209486689817606,-0.00625875293134626,-0.00250035069934862,-0.0137236331739816,-0.00492601403191495,-0.00547704689669382,0.00904394952668475
"3246",0.00222387007607705,0.00244172692033962,0.00067202971151592,0,0.00128820184693623,-0.000179126907213889,-0.0032611712703291,-0.00371294214239082,-0.00188402173913049,-0.000640183169661301
"3247",0.00775022481673382,0.00819305774095036,0.00688253560933849,0.0100302696195689,0.00293054264295867,0.000447634961338705,0.00392640327360039,0.00546592143956204,-0.00479165802266368,0
"3248",0.00226570066581577,0.0010983032437013,-0.00166712095572419,-0.00300226404089576,0.00584416888985761,0.00187942289776943,0.0120586425499201,0.004200457373154,0.00481472855537302,0.00576553466334007
"3249",0.00445757243941447,0.00153575427430774,0.0020040323543582,0.00115819048246379,-0.00290511010421401,-0.00259034505436984,0.0032202246602171,0.00196853645427653,-0.00529991268694952,-0.00509556275296941
"3250",-0.00370870940901646,-0.00569554708303066,-0.0095000853962226,-0.0157334395195967,-0.00213193605010409,-0.000806042621138037,-0.00278200245839511,-0.00294690926710228,0.00620397073950696,-0.0198463287199427
"3251",-0.00849472371349946,-0.00793126175449432,-0.00201913822928435,-0.000235087881814922,-0.0133329502301776,-0.00359033238451567,-0.0148068879826152,-0.00270929288186772,-0.000507819523372866,-0.00130635779152333
"3252",-0.00670666751570059,-0.00421947746465456,0.00387791506578727,-0.00517276307417114,0.0209675924338519,0.00891810156956652,0.00609891242904959,-0.0019759370331307,0.00957985388677685,0.000654066522213448
"3253",0.00617029394041646,0.00958964503067627,0.0112529234796681,0.00756324509713302,-0.00998536154134144,-0.00383930882488581,0.00389690869313508,0.00222725231174592,-0.00136584716148491,0.0156862734681336
"3254",0.00179808812930649,-0.0017671346984004,-0.00398602966919126,0.00445692621978799,-0.00486405153782665,-0.00233030965625303,0.000862671363753398,0.000987548869418653,0.000575885409960897,0.00193043642338497
"3255",0.00913392150769154,0.00885149537135455,0.0115057951450779,0.00583835801069088,-0.00553476275080178,-0.00305444790988507,0.00172384448168894,0.00666022259127996,-0.00992809352517998,0.00642265108196249
"3256",-0.003144069139142,-0.00438687220328426,-0.00560502629182014,-0.00394707642766878,0.00216830593544448,0.000810864874157824,0.00204335724428173,-0.000980261927361004,-0.00029060457384833,-0.00127634574400448
"3257",-0.00111515024699682,0.000440559543400498,-0.000497400021302163,0.00349648733708374,0.0000720727871488247,-0.00117039627102355,-0.00601054128132106,-0.00171687972179868,0.00283470703830924,0.00447288663458867
"3258",0.00283871673349889,0.00484482882557136,0.00215626407172631,0.0146341505319771,0.00786117860168023,0.00414667854217177,-0.00971811581308291,-0.00196563429450769,0.00688553303699702,-0.00445296900902392
"3259",0.0086189827615677,0.00832778792930711,0.00248261390356963,0.0173992263926959,-0.0164579283097778,-0.00790026894619378,-0.0130847134121639,-0.00467746464010688,-0.00352724594770004,0.00894570834782171
"3260",0.000599144402045448,0.00912847591431287,0.00264155902433205,-0.000450004420986527,0.0115678809339197,0.0058819561461454,0.000994375318600138,-0.0029680740933401,0.00447887041358164,0.00506645466891054
"3261",0.00687003104198025,0.0133553161065143,0.00459899428795008,0.00848459952967739,-0.00899033471348387,-0.0046779362080549,0.00642034156013294,0.00620199952358136,-0.0000719884917945723,0.00693133829067927
"3262",0.000219264571326372,-0.0070603800010266,-0.00215628679920121,0.00911986963188904,-0.00137888464483715,0.0000904368200618233,-0.00852802279318632,-0.0066569372801798,-0.000215750873923115,0.0043804543080963
"3263",0.0000624929395611762,-0.00107729171589399,-0.00398935448354121,0.005422537738208,-0.00821234421382788,-0.00271148138613553,0.0129580037400781,-0.000992723425900066,0.000072002016833439,0.000623031858375089
"3264",0.00409893236374703,0.0002156688673145,-0.00100127441960518,0.000449469286755155,0.001600019095229,0.000780514420526401,0.0082708398819471,0.0084471599886824,0.00258956257834675,0.00435869731147753
"3265",0.00438425921664121,0.00345048181970076,-0.000668275120421002,0.00202156754409133,0.0013190384526931,0,0.00623422730159007,0.000985467132060824,0.00100444106025099,-0.00123988358548832
"3266",0.00152775042452635,0.00236408177929248,-0.000835851964950507,0.00134492506277595,-0.0014636701121109,-0.000906650424909339,-0.00565214439720996,-0.000157303878370874,0.00308194515246707,0.000252270433905188
"3267",0.0000311265085102264,0,-0.00401536817755332,-0.00223863619067044,0.0028582763190248,0.00172439762894983,0.00273289285626821,0.00262193709928171,0.00943199019861352,0.00441361916771754
"3268",0.00532323776648513,0.00385932030248637,0.00268766473347792,0.00717971759229852,0.00241141768920072,0.0014496019922936,0.00534178161419874,0.00679919860374878,0.00785730139853325,0.00753289391086009
"3269",-0.000247786338546718,0.00384456970287328,-0.00184280502175216,0.00400981030264602,0.00109375887348762,0.00144764963979749,0.0027108855206035,0.0064933767775861,-0.000351193975586694,0.0018692213002629
"3270",-0.00551314527289282,-0.00680850429536406,-0.00889563274573513,-0.00665625961490168,-0.00364120003141988,-0.000632396451354711,0.000756921065687033,-0.00206447196973514,0.00210779874787059,-0.00186573383084565
"3271",0.00242925808725336,0.00599824262356807,0.00321766185992001,0.00223354587803759,-0.00979404371326453,-0.00361593777248559,0.00583530142226918,0.00310320730784053,0.00189293269673496,-0.0062304676779108
"3272",0.00935187127606518,0.00787912922421707,0.0104659245442775,0.0202808028745636,0.0112933462523963,0.00462700353747403,-0.0110656781181514,0.00206242247327992,0.00734781696351927,0.00125391849529799
"3273",-0.00757218177576313,-0.0107755098234247,-0.0110257312525743,-0.0185669610905006,0.01540026156853,0.00668303248024538,0.00716998997586371,-0.00205817764145821,0.0132685240695074,0.0118973074514714
"3274",0.00381507455694985,0.00363101973698132,0.00354723531942613,-0.00244831015044711,-0.00567855463214828,-0.0010766695174883,0.000862926754172655,0.00232027829556136,0.0104894967058171,0.00185649752475237
"3275",-0.00281186190530947,-0.00574595843115333,0.00168322374782659,-0.000669345469804461,-0.00491580766498134,-0.0014369164946072,-0.0101303828816522,-0.00360093716501375,0.00393515166520908,-0.000617726953815456
"3276",0.00532966906831245,0.00192636675545765,0.000168051382735124,0.00580484211486954,-0.00661079801315567,-0.00233835951775685,0.00239513395986868,-0.00722755651930396,-0.00750152052779929,-0.0148331273176762
"3277",0.00678054385093763,0.00299081391940703,0.00705641330564499,0.00665923719999384,0.00351026086771444,0.000721255729183579,0.000543133772920923,-0.00078017813394593,-0.00565165459858608,-0.00439146800501888
"3278",-0.00287768261451493,-0.00489882544544595,-0.0070069692347049,0.00529227229106888,0.00889071999789626,0.00216190795904558,0.00868421313478418,0.000520515939787414,0.00602619328922938,0
"3279",0.00687729726941355,0.00449484131646471,0.00571241441437409,0.0155735643938337,-0.00303351466374435,-0.00116841324456896,0.0106544643628426,0.00546165144821487,-0.00741948791996483,-0.00756143667296783
"3280",-0.0015246040148672,0.000639256120133824,0.000334070207346215,-0.00561554814723186,0.0051441597066777,0.00197985737543038,-0.00383348494011315,-0.000776035686098964,-0.000891544326973026,0.00444444444444447
"3281",0.00225986057170613,-0.000638847732810643,-0.00367403320403992,-0.00781932593510881,0.00663124787118186,0.002514836161426,0.00887219143884921,0.00336521119964783,0.00583424386252673,-0.0050568900126422
"3282",0.00831835190894159,0.00554016937213131,0.000670515440160502,0.00634857641216202,-0.00315044859117464,-0.00206071240251515,0.00741692983440045,0.0064499262945148,-0.00156950328228833,-0.00127064803049548
"3283",0.00311267389171355,0.00487391095977574,0.000669998617085277,0.0056558378504179,-0.0085481647695157,-0.000807905694298561,0.00115689468581448,0.00410150373710394,0.00184542412474098,0.00318066157760799
"3284",-0.00195823342305934,-0.00801348128755508,-0.00535656887638147,-0.0253082295422152,0.0105055218237569,0.00395322957267874,0.0101901670606306,-0.00663774191197808,0.00109157455189557,-0.00570703868103994
"3285",0.000120720929629892,0.00063776125118209,0.00454388663352967,0.00821121668140612,0.00351353474882377,0.000179056461237614,-0.00571964464551156,0.00411215051067537,0.000340656932647843,-0.0133928571428571
"3286",0.00114688642773109,-0.00403650135268774,0.00117274476327234,-0.0103455941509641,0.00700168623913511,0.00250538539225453,0.00596167120324864,0.00204764183152695,0.00224812327635981,-0.0084033613445379
"3287",-0.00889313509130618,-0.00234643169898918,-0.0038486917843138,-0.00800709001129607,0.00808851611927275,0.00357010918322431,-0.00228740138394179,0.00229894228327554,0.00584557523944995,-0.0149934810951761
"3288",-0.0160293319332613,-0.0205259590025008,-0.0179741526220804,-0.0345290563193338,0.0155546874731036,0.00675914047185922,-0.00479364181141428,-0.0127422635106216,0.00682530765847567,-0.0185307743216413
"3289",0.0104791418454446,0.00873165438198131,0.00889498922348486,0.00836030421661405,-0.007831361575109,-0.00335677817984192,0.00429320142408396,0.00129067774754521,-0.00892678002125047,0.00472016183411994
"3290",-0.000826043276320521,0.0012984108822276,-0.0032214122583295,0.00483658399892262,0.0097790052222031,0.00478621535374724,-0.00312789096219601,0.00567150276215589,0.00541787199193089,-0.00469798657718123
"3291",0.00324539213698727,-0.00129672719752316,-0.00136080740599354,-0.0148981134834871,0.00013868184933119,0.000970434479244942,0.00125508642285377,-0.000256269854291502,0.0000673177928653956,-0.00876601483479433
"3292",-0.0181579409958159,-0.0157974309889632,-0.0163515801850939,-0.0202419232999226,0.00912970707062066,0.00502338600872831,-0.0121174184516289,-0.00410255509830115,0.0057924226726449,-0.00816326530612244
"3293",0.00742863494221568,0.000879567893601552,0.00761903388901453,0.0111612520740343,-0.000810158628212987,-0.000851665898069953,0.00306644525517741,-0.00102993664695727,-0.00649568731673889,-0.0185185185185185
"3294",0.0152411011355513,0.0158172190162569,0.0151229155854107,0.0258337162767477,-0.0134668971058823,-0.00580031554842142,0.0102256174753554,0.0048970176752936,-0.0130089511120994,0.00139762403913335
"3295",0.0115480752854902,0.0114619088852357,0.00897236787122901,0.00572347069933188,-0.0109349348304075,-0.00433114808796309,0.000208643952275045,0.00051282892436344,0.00122931099231849,0.0153524075366365
"3296",0.00336487782430317,0.00171044246794572,0.00755033471921118,0.000910510871284131,0.0045069585409605,0.000710166635423004,0.00375598119378706,-0.000512566065659414,0.0053883977533018,0.00412371134020617
"3297",-0.00532967646223181,-0.008751324999831,-0.00965859211977571,-0.0138730713250126,0.0124779871185379,0.00479070753451727,-0.000415809771089681,-0.00461664699596231,0.00264585492452607,-0.00547570157426425
"3298",0.00746539097591192,0.0025840478828647,-0.00117701531755454,0.00553499735918916,0.00276953045381489,0.00194241193563549,0.0100863268384814,0.00566868613223792,0.00257124986804746,-0.00894700619408118
"3299",0.00173294652095879,0.0060136801552948,0.00505050410780439,0.0130733995747947,-0.00504041567981228,-0.00237934693005615,0.00813264183186679,0.00358688754167891,-0.00344195185856722,0.0034722222222221
"3300",0.0064428080399217,0.00576435966343181,-0.00485767569065076,0.0135839551834362,-0.00506595017450495,-0.00256171174115027,0.00796475223596937,0.000510682356676728,-0.000812752246708404,0.013840830449827
"3301",-0.00106695939809442,-0.00785397690223211,-0.00875268544621122,-0.0131784800834763,0.00383633517902138,0.000885620955479283,0.00678762087947393,0.000255223964669593,0.00569345289314205,0.000682593856655256
"3302",0.00160214551515936,0.000855770161738434,-0.00747154323348964,0.000452724825878104,0.00437729186691893,0.00247759618246035,0.00905608984443496,0.00867343342949622,0.00417842687092507,-0.000682128240109159
"3303",-0.00257702825816741,-0.00448907627735451,-0.0148845448118777,-0.00656115255645673,0.00684884444735423,0.00158868020474645,-0.000697970664390146,-0.0035406226365815,0.0128188187919462,0.00750853242320826
"3304",0.00478117978676074,0.0057976926925265,-0.00173670217705524,0.00728761108863663,-0.000068652314647033,-0.000176278483056347,-0.0125736347311632,-0.00304581523019831,0.00583121712726231,0.00948509485094862
"3305",-0.00410810076505885,-0.00597773198707041,-0.00643705783027193,-0.0156001910728693,0.00783352910720003,0.00290856200218603,0.010813515224104,-0.00381877636813255,0.00408466320964895,-0.00402684563758393
"3306",-0.0102983298730508,-0.00279213024142766,-0.00840479981402165,-0.00574185072685018,0.00934052528582319,0.00404247470302055,0.00189968666446183,-0.0020445021867882,0.0150252144865768,-0.00404312668463613
"3307",-0.0331654364772118,-0.0432910215776544,-0.0337277014263615,-0.0374220915704251,0.0149284576648472,0.00778995160816343,-0.0133718959600075,-0.0197183324066023,0.00898512622466319,-0.0189445196211095
"3308",-0.0303021852536747,-0.0229626008158278,-0.00164472917725533,-0.00791931086011777,0.00532460375242128,0.00277911928604002,-0.0268028695497853,-0.0107104156142139,-0.0178742588986933,-0.0186206896551724
"3309",-0.00367813132197181,0.000921628994235091,0.00494237165425981,0.00798252697266366,-0.00529640250775421,-0.000519566050983244,-0.0104967559124817,-0.0105624948312235,0.00437050219757662,-0.00983836964160234
"3310",-0.0449116597365058,-0.0303867778650727,-0.0342441068723104,-0.0239980989444386,0.0108487081535571,0.00485266487176705,-0.0524104823069581,-0.0240192967046704,0.000194836655226238,-0.0170333569907736
"3311",-0.00420159335836701,-0.00807209288418276,-0.00113167483122412,-0.00368815598952044,0.0225835223048778,0.0112108284095724,-0.0312568791560756,-0.0213287903680033,-0.0364934740259739,-0.0173285198555957
"3312",0.0433064030565811,0.0179511760230457,0.0126510959006805,0.0217176822931475,-0.00735739563819504,-0.000683165246036954,0.0481692243227316,0.00558810451230629,0.00552629715843445,0.0227773695811904
"3313",-0.028632345988727,-0.00893485234892677,-0.0128659982779956,-0.00676338807140464,0.0155256850294621,0.011620030203247,0.000109172198041296,0.0133370084178119,0.0314343303907707,0.00215517241379315
"3314",0.0420329868267011,0.0360616145976007,0.0217227082900311,0.0177528997167657,-0.0106186893934238,-0.00219597186577214,0.0382012211576799,0.0235811182574088,0.00175453246965063,0.000716845878136363
"3315",-0.0332416318186808,-0.031600575982304,-0.0181179278773111,-0.0210273969014174,0.0248916957411707,0.00888783595461895,-0.0217618575872334,-0.003750426128449,0.0216009400207333,-0.0107449856733525
"3316",-0.0165311137369377,-0.015133587127014,-0.00960271735351292,-0.0205028255014883,0.0520440108834674,0.0101519452540602,-0.016980220658078,-0.0188221709390026,0.000380963858627181,-0.0325850832729907
"3317",-0.0780945080475549,-0.0871548959048142,-0.0509505915882864,-0.0682781074044917,0.0271030241629875,0.00896992161905974,-0.0741226279124959,-0.0570019851747433,0.00165023798825326,-0.0778443113772455
"3318",0.0517449477200351,0.0360336318441716,0.0298477980785015,0.0508157987082745,-0.0512580480367424,-0.0183568926153396,0.0386113152031951,0.00610286167445473,-0.0211013373183111,0.0316558441558441
"3319",-0.0487483626877869,-0.0558517218920352,-0.0338456002982125,-0.046576833265209,-0.0367976980975238,-0.00997910349587405,-0.0582082150347392,-0.0283073450178859,-0.00356035094666884,-0.0180959874114871
"3320",-0.0956772613785927,-0.113471359822084,-0.0980471007715304,-0.100106782587216,0.00619690933897465,0.000508300828530261,-0.0974167603071193,-0.103448270592329,-0.039888262711738,-0.0400641025641025
"3321",0.0854862319939624,0.0606612905043435,0.0328125133233683,0.0720854416965411,-0.0226032304067226,-0.0065187560307709,0.0853284308911568,-0.0135941920931343,-0.0305162339374359,0.0108514190317195
"3322",-0.109423655124521,-0.113239960662234,-0.0659174018185277,-0.124792455870564,0.0647656371007326,0.0264166262802079,-0.168699954026307,-0.0988234920045739,-0.011446119566207,-0.060280759702725
"3323",0.0539920099937139,0.0451467253883813,0.0490512730224493,0.0689220041521224,-0.0666830199129139,-0.0250727204319019,0.0469907659925841,-0.0193957337079046,0.013555485834196,-0.0158172231985941
"3324",-0.0506329333339818,-0.0688059397979771,-0.0211732745069986,-0.0863650588904465,-0.0564126019976608,-0.0138804817850782,-0.0984000266495013,-0.0928109729441079,-0.0199219910827807,-0.0330357142857142
"3325",0.00212496810922769,0.0218687965462918,0.0139701966292072,0.00776948874572714,0.0272254815296109,0.00328150171078478,0.000471100862792673,-0.0612159433256795,-0.0189055014692003,0.0212373037857803
"3326",-0.0430941701749346,-0.01264590472113,0.0024444680077409,0.00738843034004999,0.0751955682963028,0.0254776385272615,-0.0437922955947413,0.0236713647440396,0.0149957121484352,-0.0108499095840869
"3327",-0.0255681792137884,-0.008210170851641,-0.0104190069628446,-0.0239158343674666,0.0412091908266699,0.0118349221064422,-0.0505580117811998,0.00334731273147448,0.0441795871516695,0.0118829981718465
"3328",0.0906032647670119,0.0894039600785337,0.0694445109276576,0.0751388490113072,-0.0186144803395161,-0.00680221298569028,0.0800484020912082,0.0930640970784973,0.0485303544388853,0.0216802168021681
"3329",0.0149701833313418,0.0407294644454257,0.0188521120706182,0.0352476684856273,-0.00227112815592379,0.000584645359708924,0.0549027246964815,0.0650602512143974,-0.0136896419956835,0.0167992926613616
"3330",0.0583897595012151,0.0487733807637045,0.0328947169377323,0.0378632132018168,0.00492192525237822,0.002420667772979,0.0741536122733066,0.0282806118894561,0.012822220499229,-0.00347826086956515
"3331",-0.0297856485828085,-0.0345308871970851,-0.00119427534282046,-0.0568440105146153,0.0266928095174155,0.00741122061234334,0.00128357948382396,-0.0352036366302383,-0.00646048660726684,-0.00349040139616064
"3332",0.0324757222262593,0.0187482532395389,0.0121562302676208,0.01649193150483,-0.00822902297877626,0.00231429367901903,0.019943026437049,0.00836199565726536,0.00440064367816095,-0.00262697022767067
"3333",-0.0149053477718435,0.0002831953295932,-0.0275644704246693,0.00678462520710532,-0.00811687629248781,0.00181431191762105,-0.0283518497883229,0.00904629620280839,-0.0318466849574507,-0.0122914837576822
"3334",-0.0450048979336971,-0.0467025093888636,-0.0475804605704716,-0.042777684440564,0.0140107048864517,0.00407133799049508,-0.0659767569063738,-0.0362346586816086,0.00945622405694913,-0.0284444444444445
"3335",0.0230754255165595,0.0190023573042193,0.0127550996903834,0.0336700549201294,0.00634587529037112,0.000164053610447468,0.00430911901207187,-0.0104650852944225,0.0163934228784226,0.019213174748399
"3336",-0.0144541988287852,-0.0203963583765886,-0.0224601444923543,-0.0189517032637314,0.00237937513967679,0.000738833243623116,-0.0156298978346084,-0.0336857722805298,0.00493745904953746,0.0251346499102334
"3337",0.0671662219954399,0.0475908003136436,0.0590508748002796,0.0546332159856917,-0.00261131898099176,-0.00451053027387638,0.0750311064467535,0.0381029516962397,0.0277105218883926,0.00525394045534155
"3338",0.00101947017773707,0.00454292669478429,0.0107461229525387,0.00515169968206397,-0.0104723479267606,-0.00444838254916524,0.00970173181356415,0.0394376513755572,-0.00535448733571875,0.00696864111498252
"3339",0.0335683431612204,0.0146975764625425,-0.00240717690656544,0.0102505341176606,-0.00727594213142158,-0.00124142273913286,0.071561682488946,0.0202855150895977,-0.00890796630579194,-0.00259515570934266
"3340",0.0152173714965285,0.0239553413878955,0.0130705722980813,-0.00366403459052778,0.00181706632503831,0.00215430314225507,0.0556745023835563,0.0261414303111067,0.0261235574312406,0.0026019080659152
"3341",-0.00913015879142376,-0.0141457085925093,-0.00416832813663603,0.00141449661856963,-0.00912992892203224,-0.00214967209690198,-0.0406946208037019,-0.00717616525115194,0.0171403488923014,0.0173010380622838
"3342",0.0294929467621732,0.0187636316379094,0.0183376587307822,0.0228812619783516,-0.000244013621497174,0.00132563154438836,0.0264305233709998,0.00542098010660719,0.00786809347950945,-0.00850340136054417
"3343",-0.0212481029475734,-0.0392739759094489,-0.00998231150838602,-0.0256834580933755,0.0264891055066152,0.00893617101560396,-0.0378523476211189,-0.0287562888330475,-0.00510196112437744,-0.0205831903945112
"3344",0.00482425802820696,0.00281920625756293,-0.00850143253194413,0.00538548954046902,0.0113568991408131,0.00106597541124342,-0.0112406055551213,-0.0074019146513068,-0.000864992244733132,-0.00262697022767067
"3345",0.0270153530438513,0.0334551593858361,0.0133598803951214,0.022272324237756,-0.0134046514552736,-0.00262139226526104,0.0297739107837502,0.0294556039319709,-0.0194174748876239,0.00438981562774354
"3346",-0.01761797031896,-0.0136017254993893,-0.0153482503053757,-0.0126862013663323,0.00804490807177194,0.00262828202342802,-0.0362727217273517,-0.0130387516830515,0.00712612694782822,-0.0166083916083916
"3347",-0.0303632095612731,-0.0206839532440098,-0.00939251392664298,-0.0276534673841202,0.0125915793830718,0.00278531259978099,-0.0182735868497295,-0.0264219386860173,-0.00682527251393739,-0.0471111111111111
"3348",0.0221945689385128,0.0152069310627412,0.0173492019862005,0.0272908711650941,-0.0102166155279998,-0.00310439136338736,0.0159744905142423,0.00980013182525785,0.0196708592165005,0.0139925373134326
"3349",-0.0000717818086514166,-0.00776693456136479,0.0013881050999287,-0.00363523274802269,0.00530857631484483,0.000655657574721413,-0.00916052150005198,0.00373271221196769,0.00995486328955342,-0.00275988960441576
"3350",0.0139387609195352,0.0123007783890858,0.0077227428958202,-0.00140335233329325,0.00234670848110197,0.000245586066749182,0.00413957708282031,-0.000371833849167391,-0.00428552110409031,-0.0129151291512916
"3351",0.0144184910535579,0.0143606822941515,0.0137551626250407,0.0202359886775731,-0.0186138090042597,-0.00532172622199012,0.0316065441133615,0.0171131065150638,-0.00664043904722345,-0.0186915887850466
"3352",-0.00459854802880921,0.00707879663351374,0.0145376792194676,0.00192836964071885,0.0115113297454743,0.00436246892131886,0.00905809612130026,0.00658377728160797,-0.00445656108512704,0.000952380952381038
"3353",0.026178579886365,0.0267638627434987,0.017577346690028,0.0291449267118005,-0.00518897597504242,-0.000491657942069956,0.015313563932623,0.0243458804204391,0.00553344952831258,0.0180780209324451
"3354",-0.00931067050279188,-0.0184307270035744,-0.0281637220662144,-0.0211060477040499,-0.011676709110597,-0.00237786843496368,-0.0111817978959757,-0.00638525989898464,-0.0181165712759925,0.0186915887850467
"3355",-0.0264734602432194,-0.0206545609110421,-0.0175811560578513,-0.03602622343947,0.00856310842595809,0.0013822749612038,-0.033925132704249,-0.0199928483209154,0.00617125932925822,-0.0128440366972478
"3356",0.00275827204090495,-0.00109544374983017,-0.00491642696561245,0.0107588952064777,-0.00470362005877267,0.000164364139649376,-0.00299443640685049,-0.00546446445131643,0.00350480037241718,0.0120817843866172
"3357",0.00923931665982503,-0.00219370652040352,0.0096838519972684,0.00560220546217072,-0.0064010594080981,-0.00073940991628163,0.00477819286845205,0.00366294285011515,0.00424103790048735,0.0257116620752984
"3358",-0.00677870494884525,-0.00741958132599008,-0.007633559021617,-0.00306402656752314,-0.0161357855809483,-0.00369939752058501,-0.0165761915449618,-0.0113137855469899,-0.0128555890484265,-0.0196956132497762
"3359",0.0120667690657279,0.0166113157015229,0.0149900704423751,0.00810279180220941,0.0167062646423475,0.00610611837023489,0.0132634161328704,0.0184569515255051,0.0153507520984728,0.00639269406392695
"3360",0.0165462542525854,0.0166121764765872,0.017100688820046,0.021064308227752,-0.013000957569097,-0.00328059431042038,0.0238613836229253,0.0224718918619804,-0.00601029187688384,0.0208711433756805
"3361",0.00020510148946129,-0.0048218242444994,0.00955293469599394,-0.0065146987999174,-0.00780592293519777,-0.00279764359489143,-0.0141163495660102,0.00248151455427492,-0.00623363678136934,-0.0133333333333334
"3362",-0.0199315050681369,-0.0123823350200855,-0.0130582795686577,-0.0038252088283165,0.0102643635592363,0.00330055976788213,-0.0459272896529588,-0.0275814238776146,0.00388906666527511,-0.00810810810810814
"3363",-0.0176859050894581,-0.0136276766684582,0.00479386952469163,-0.00191987965241502,0.00699629443803462,0.0020561338419951,-0.0236443574788023,-0.0152727923759035,0.00962265100823889,-0.0099909173478655
"3364",0.0119673303210499,-0.00828955125068231,-0.0148855360195997,0.00384725591902502,0.00978735299669387,0.00155935677107633,0.00464037082080693,-0.00443126395712379,0.00885006177930348,0.0174311926605504
"3365",0.00459701600979745,0.0016717910270807,0.00174350223676001,-0.0136873907725067,-0.00257265184610778,-0.000655535187989109,-0.00461893723921891,-0.00964390060318909,0.00564381343610254,0.00991884580703339
"3366",0.0304596005916291,0.0445062188204637,0.0249468665265471,0.0391339704865852,-0.0219542274440506,-0.00615005221966791,0.0582946694509008,0.033333321889516,-0.00756414965502994,0.0285714285714287
"3367",-0.0102711969626738,-0.0143808570434319,-0.0116980631014117,-0.00801275757095932,0.00374122380809672,0.00280531887916369,-0.0112358395179575,-0.00144982090979595,0.00965021194111237,-0.00260416666666663
"3368",0.0169880442044297,0.0224264980534858,0.0150819916545704,0.013193368843696,0.00299390246664988,0.000246734181868158,0.00970051227268254,0.00725959274279542,0.0023742786550065,0.0174064403829417
"3369",-0.00690393747770979,-0.00845665158740994,-0.0107202880622216,-0.0114270946278935,0.00249772972055085,0.00065813943786952,-0.00137236654096085,-0.0100901205235654,-0.014576338217176,-0.0042771599657826
"3370",0.00189909283510747,-0.00266530673369203,0.00133076249699848,-0.0206988698054134,0.00601608110696228,0.00189060842110389,0.013606271920801,-0.00327632861658333,0.00591683821263467,-0.00773195876288657
"3371",0.0123204526819634,0.0253875128402588,0.03398522998176,0.0219598675808801,-0.01340983470375,-0.00262554073393473,0.036474619549415,0.0365229995509746,-0.0142148636756079,0.0103896103896104
"3372",0.0148790792866915,0.0138129461020329,0.0128534745287201,0.00322313292248255,-0.00183670959993176,0.000822694497789156,0.0192308148376461,0.00845670620548811,0.00180243645846501,-0.012853470437018
"3373",-0.00184497583633136,0.00925435295810217,0.0130529493666196,-0.00696104081879789,-0.00368046210434048,-0.000904143344512387,0.00410719860636743,-0.0027952514852676,0.00335034137890799,0.00520833333333348
"3374",0.00445595214652239,0.000509446485465137,-0.00841090541624345,0.0172552702109701,0.00714158721870572,0.00320860139132106,-0.0103540947515436,0.00875970429676975,0.00735841573486007,0.0172711571675301
"3375",0.00404169032652724,0.0224033037468216,0.0151597088697628,0.0230585164179555,-0.00673267499427832,-0.000394212082825418,0.0231206867953475,0.019451150029032,0.00460376883914382,0.00594227504244493
"3376",0.00828007719103896,0.0114542012321317,0.00444443186142518,0.0238342835950285,-0.00363574063423533,-0.00164241467466464,0.0089635409746458,0.0252129514573673,-0.00647682985514275,0.0109704641350212
"3377",0.0133083461235106,0.0295420327686855,0.00690264682839925,0.0232793331388748,-0.0132970160698368,-0.00592247432059911,0.0300300135525986,0.0312396095852701,-0.0184501838210265,0
"3378",-0.00262675337908724,-0.00310850183458411,-0.0112497599973835,-0.0140949604159364,-0.0144791812699764,-0.00397185592007787,-0.0085033542843701,-0.00902352005641893,0.0105262715341001,0.00834724540901499
"3379",0.025629500793557,0.0191892849070205,0.0144000767787158,0.026335570795549,-0.00712319871697242,-0.00498467638116507,0.036387971548909,0.0198373600063886,-0.02027532254635,0.0198675496688743
"3380",0.0120875046654561,0.0115320293497685,0.0147213179967907,0.00610948678742806,0.00384337943109836,0.00108549819259829,0.026362515667872,0.0191325954796409,0.0108221381818283,-0.00649350649350655
"3381",-0.00745664427818782,-0.0155885456661125,-0.00518141579093911,-0.00680107510660422,0.0113584961881372,0.00358635381150507,-0.0161253216862736,-0.0134542038069074,0.00964183565212973,0.00326797385620914
"3382",-0.00557998368777679,-0.00354531908457989,-0.00052080177154501,0.00733669906076417,0.0148274399494048,0.00747942457205952,-0.0255209273176124,-0.007294757617751,0.014324767900433,0.00651465798045603
"3383",-0.0576489707513297,-0.0600094501369361,-0.0420357316955461,-0.0521970138927943,0.0189007997795123,0.00354694210810047,-0.0631906378782332,-0.0578274572836955,-0.0072140854038113,-0.0323624595469254
"3384",0.0119756803463431,0.0181679735531781,0.0179509584773114,0.021260195437363,-0.00964118662957103,-0.00221935373554327,0.035778216505258,0.0267887890148186,0.00141631874756021,0.00418060200668879
"3385",0.00933565772188905,0.00963476037823074,-0.0109159758309445,-0.00908173584969074,0.000554414933942038,-0.00082377387929744,0.0115034973281549,-0.00825630592771898,-0.00178325549696379,0.00915903413821817
"3386",0.0192477141878538,0.0119284039797019,0.0192412779088764,0.00636456228015692,-0.0153333889325676,-0.00206110781085989,0.019714145968118,0.0116550220907274,-0.000492835575767514,0.00825082508250841
"3387",-0.00415391792027364,0.00319246062886869,0.00445235959207979,0.00961297772863601,0.00412753881257322,0.00156973253351733,-0.0135331267359053,0.00592489935526097,0.00191061941448378,-0.0049099836333879
"3388",0.000385002948950941,-0.00758866622221144,-0.00177310277400344,0.00050112753695819,0.0105879772268502,0.00222710162048223,-0.010656522812962,-0.00589000168805687,-0.00196846090020264,0.00575657894736836
"3389",-0.00571488387496744,-0.00370009857671172,-0.00479573720773963,-0.000250488354620604,0.000801120721800386,0.000329272278315473,-0.0126283981247163,-0.01547066925223,0.0110330001530756,0.00817661488143906
"3390",0.00641524512125113,0.0143600399693002,0.0067820989966465,0.0122745998133567,0.000123327974909326,-0.00090506255619216,-0.00188095619465689,0.00752692060578486,0.00646221426850113,0.0105433901054339
"3391",0.00460365509630378,0.00585789587849894,0.00265912072327601,0.00965105171987135,-0.00683453859685279,-0.000329470332892989,-0.00301500926028264,-0.00435514477014409,0.00841965009194134,-0.00481540930979141
"3392",-0.025508699648112,-0.0266925024676659,-0.0208628001969094,-0.0132353189518459,0.0107252540869172,0.00189478562547052,-0.0286039431220005,-0.0211978679724223,-0.00348391406736948,-0.025
"3393",0.0107205322028541,0.0157068308225672,0.0113758936190702,0.00422260328974677,0.00288299843358897,0.000164436597315687,0.0123233869468826,0.00446892674177124,-0.00060271852692162,0.00909842845326714
"3394",-0.0237514526070287,-0.0179186049131759,-0.00964108229391469,-0.0121197378184517,0.0107032453948561,0.00271291435958632,-0.0198617202507195,-0.0102669588847596,0.00446314829077532,-0.012295081967213
"3395",0.0146974757705778,0.0119971013245237,0.000180259596533894,0.00450676025304864,-0.00314668987254219,0.00098382953433318,0.0186952461498193,0.00242046883942448,0.000540482789620489,0.0165975103734439
"3396",0.0128095961559194,-0.00222277094478773,-0.010093763518385,-0.00324020446760243,-0.004856507211772,-0.00180192154496317,0.0114219859685722,-0.00586407271135569,0.00444091686848336,0.00489795918367353
"3397",0.00700483221867909,0.00816826692236283,-0.00200285877650619,0.0112527376217686,-0.00194214388198055,-0.00156048132695796,0.0224591933239477,0.0156141323850161,-0.00448108993490737,0.00812347684809089
"3398",0.00550690393987163,0.00932975693591942,0.00656808964480771,0.0227498027386202,0.00104034099575334,0.0012338791927049,-0.00310255714473595,0.0143492235632483,0.00216061103590848,0.00402900886381952
"3399",0.015437332571179,0.0184869370351026,0.0128693678763592,0.0430367010871204,-0.00409562052881696,-0.00147881881374479,0.000124402352400299,0.00707298211016538,0.00598874131006677,0.00802568218298561
"3400",-0.010313816430808,-0.0157630765646781,-0.00894774500809337,-0.0166898705769558,0.0140560176794908,0.00320878544484571,-0.0190440405686808,-0.0170568374208426,0.00631025732373525,0.000796178343948961
"3401",0.00764860956357905,0.0111623152429583,-0.000722300456440839,0.0259312129151916,-0.0039949165325166,-0.00155824002168115,-0.00101503907931721,0.00510387204307716,0.00621156556720881,0.0127287191726333
"3402",-0.00569293969729834,-0.0139188391609714,-0.00487893024936759,0,0.0159221139099186,0.00320351391736651,-0.0055887260025832,-0.0135410306842894,-0.00270439773542008,-0.0117831893165751
"3403",0.0102105839914772,0.0109515940618155,0.0130742872707463,-0.00643377757352959,-0.00502481965422197,-0.00196506263555152,0.00281006769971381,0.0061770874471303,-0.00259389840848034,0.00635930047694755
"3404",-0.00865898910452056,-0.00481466045222279,-0.00519808200039285,-0.00670677582299828,0.00330675792975166,0.00106652658742679,-0.012355079777307,-0.00920873072510819,0.00124116081043613,-0.0102685624012638
"3405",0.0129590212140345,0.0164489598451862,0.00792790990990988,0.00139690334349485,0.00143811803142824,-0.0000819076418656639,0.00760894490904418,0.0103270410843739,0.00466356569056314,0.00478850758180371
"3406",0.00918721257613631,0.0128510471204188,0.0126922240381162,0.00302257628563485,-0.00466724362418725,-0.000327920082654809,0.0103674114142491,0.00306642783482847,0.000881332617882036,0.0119142176330422
"3407",-0.00329340122625077,-0.00469924800988619,-0.0102383403269782,-0.0141400095999077,0.00474926110929319,0.000737865138610294,-0.0108944032039501,-0.012228282939188,-0.00945168508751182,-0.00784929356357922
"3408",0.00289902053674718,0.00660996207247511,0.00160513643659699,0.0056430991216343,-0.00209415633635968,-0.000245708055866656,0.0125511984243334,0.00412662438045808,0.0082380076628461,0.00158227848101267
"3409",0.0080816469029763,0.00633210615225366,0.000712268518518577,0.0128594809445872,0.00245836221412765,0.000655535718534495,-0.0118897102609898,0.00102727813342107,0.00482016825829334,-0.000789889415481859
"3410",0.00212755005854048,0.00302962013516672,0.000533790026089109,0.00923363342566952,0.000598036837167637,0.00106460510724204,0.00256013342489392,0.00547384999707834,0.0120510002100036,0.0142292490118576
"3411",0.00569202705016947,0.00302037632387608,-0.002667579583852,-0.00434588279172288,0.00298885233434754,0.000327237565509231,0.0153217294191863,0.00544408441028921,0.0152023410404625,0.00623538581449723
"3412",-0.0119317430430642,-0.00833905528557122,-0.0033880704925795,-0.00804040909810255,0.0116812610552355,0.000981383357797627,-0.00515587969600539,-0.00913705514434771,0.00882530294296791,-0.00232378001549183
"3413",-0.00644036116093327,-0.00700777839271705,-0.00107348364776327,-0.000926377952755852,-0.000058918319754353,-0.000490239233194578,-0.00758436236338622,-0.00102464368324284,0.00857886928576646,0.00155279503105588
"3414",0.00729240701443268,0.00988007574124095,0.0198817295403284,0.015530876576979,-0.00371153553695525,-0.00155302603362995,0.0115908242590592,0.00649576722463752,0.0197537720160119,0.00930232558139532
"3415",-0.00634237481191835,-0.00372699743768923,-0.00614680376092025,-0.00821730179828117,0.00691861898038182,0.00237416294005266,0.017879603053603,-0.000339703083125031,0.00834112952513033,-0.0053763440860215
"3416",0.0122987283083531,0.0114565817161563,0.000530111327089466,0.0161104944508517,-0.00170308347208503,0.00130674664395869,0.0223899948273034,0.0190282259851782,0.00751023129251704,0.00540540540540535
"3417",-0.00356788244023998,-0.014794244789378,-0.0150123457261099,-0.0126840764356023,0.00658852668449206,0.0013865614355546,-0.00508164327849181,-0.0103367583990788,-0.00740025907739816,-0.0115207373271889
"3418",0.00790215365550329,-0.0213514786802317,-0.025820297651067,-0.00688228951594416,-0.000642874221081113,0.000244482872673313,-0.00206746723952111,-0.00707550136036739,0.00908793015585352,0.00543900543900544
"3419",0.00695221367418197,0.0191800292299216,0.0204306452998106,0.00692998366990127,-0.00503480116760047,-0.000489082750897873,-0.0130391808783741,0,0.00113253523123413,0.0100463678516229
"3420",0.00386260649785664,0.00282293591262928,0.0111832974600161,0.0133057582014222,0.00953225598945884,0.00342463434013607,0.0125941938822767,0.0115371546064917,0.0212777258202852,0.00535577658760533
"3421",0.00621093828530417,0.00492608480117096,-0.000713539052558998,0.0108671954207469,-0.00874277808313861,-0.00333167497322684,-0.0037800847354027,0.0110701139480471,0.00928324298292615,0.00837138508371371
"3422",0.00668453909538047,0.00210084033613445,-0.000714030703320323,0.00313547578340523,0.00558594031474779,0.0011414707332289,0.000122414806110749,-0.00464498733666063,0.0132740680447117,0.00754716981132075
"3423",0.000717949391551453,-0.00605641742371299,0.000357270453733571,-0.0205403433681548,-0.00666591182911203,-0.0021174956243255,0.0135846319111912,-0.00200000363190678,-0.0158853010257635,-0.0134831460674157
"3424",0.00298887799917846,0.00257794715621973,0.00482142857142853,0.00250743110342899,-0.00447381989582263,-0.00106090054070906,0.00241484689151328,0.00334006436572887,-0.00345895921030315,0.00531511009870922
"3425",-0.00825465930880132,0.00467510529862336,0.00817487115692184,-0.00272849022282851,-0.011884987133276,-0.00343140645076456,-0.0144543221454496,-0.000998687000471676,-0.0536944113708465,-0.0158610271903324
"3426",0.0139423706020392,0.0223359469520708,0.0211528291909044,0.0134518920781603,-0.00909587125076938,-0.00295126008741053,0.00965536872696604,0.0103298692791276,-0.00466820045939531,0.0107444359171145
"3427",-0.0018078390331937,-0.0059171371396709,-0.00120833764888661,-0.00292465685208876,-0.0106889740529249,-0.00205563263955111,-0.0113788706804967,-0.0042875678765647,0.0236180673271447,0.00531511009870922
"3428",0.0000297448160662128,-0.0107600961538461,-0.000172882817613407,-0.00180500902527081,-0.0039067520219157,0.000494384563117345,0.000122558329554545,-0.00364366947016281,-0.00430921830241404,0
"3429",0.0031765856964765,0.00786854912910306,0.00414869504403437,0.0126581594639168,0.00251252362943144,0.00164701335556661,0.00783541855678438,0.00698144624406805,0.0216939144946717,0.0166163141993958
"3430",0.00216040549039498,-0.000459242260832271,0.00344295059390598,-0.00111604913205465,0.00715206426058934,0.00172653193981231,-0.00473762138604228,-0.000330137001859798,0.00900800536193036,0.00222882615156017
"3431",-0.00416374217907101,-0.00321617282830611,-0.00531825346854942,-0.0122904804469274,-0.00625152450327593,-0.00131317196050107,-0.0179421018766478,-0.0142007791234133,-0.0315654597776502,-0.00296515937731656
"3432",0.00311357917991262,-0.00276559121377251,-0.00362193859951698,-0.00316742074281851,0.00903928379262475,0.00287640093338126,0.00907285048763251,0.0130652653216625,0.00691393198765544,-0.00148698884758358
"3433",0.00354737328420285,-0.00924430321238745,-0.00276958629046231,0.00499314559706887,0.00599233115701803,0.000737525006636819,0.00147793243163563,0.0056216756353944,-0.00801090463215259,-0.00967982129560674
"3434",0.0101331899471528,0.0158619084642386,0.0111091648826738,0.0110659668262414,-0.00162457077169131,-0.00139213164056584,0.00787107404447318,0.00361730975409325,-0.00565840249221783,0.00526315789473664
"3435",0.00349928625236418,0.00229628019050021,-0.00137342489270387,0.0100513960241233,-0.00765375179237837,-0.00237794196155783,0.00244056956108807,-0.00229360959694436,0.00121547513812148,0.0082273747195214
"3436",0.0100255848038739,0.00801828141955174,0.00275062756577715,0.00265367088337753,-0.00382605873906816,-0.000410983133528275,-0.00937309430182209,0.00591127445966766,0.0118088510550225,0.00222551928783377
"3437",0.00218657559608393,-0.0129545454545454,-0.00925768869337606,-0.0083811424790472,-0.0170090712300059,-0.00353595422916853,0.0142541249550452,-0.0111001613587999,-0.0115619327467172,-0.00370096225018501
"3438",0.0064593857553259,0.00736817867833306,0.00536419786530207,0.0131227760925883,-0.000744284321043898,0.00165041130340304,0.00617883903616478,0.0158467759300682,0.0173802356714787,0.00668647845468051
"3439",-0.0036225298069299,-0.00937142857142848,-0.00137690194068507,-0.0221733923638506,0.00664107083786103,0.00107108385162547,-0.00963279401238737,-0.00682479269209402,0.00238626282545851,-0.000738007380073902
"3440",0.00941857742703722,-0.00115364559298581,0.00275766976904501,0.017063268588611,0.0114377585798699,0.00327778313329619,0.0010941948033214,-0.00163613409122609,0.00119028836021973,0.00147710487444619
"3441",0.0144640265866818,0.0159389924708018,0.00996902715709869,-0.00264898460593788,0.00952030385987834,0.00139548514201282,0.0182171647408234,0.0114716748243153,-0.0131316290764936,-0.0132743362831859
"3442",-0.0344143289881788,-0.0238744884038199,-0.0175288978056127,-0.0190349712262062,0.00284125864878804,0.0013116157277091,-0.0124044761962303,-0.0123137183262474,-0.00810423853094511,-0.00896860986547088
"3443",-0.00816473940824658,0.00232935010482183,0.00554302788844629,0.000451263537906144,-0.0189884502922928,-0.00556693400627206,-0.00458945313982262,-0.00492125225186135,0.00276029591895943,-0.00904977375565608
"3444",-0.0273229169246684,-0.0141761797391629,-0.00826871676604157,-0.0173658096526839,0.00614477061125807,0.00214046264805745,-0.0124969427142561,-0.00527529236653279,-0.00192692139356365,-0.0243531202435312
"3445",0.0197474176548633,0.0238095720796592,0.00347403161368764,0.0149185448703237,-0.00268719913621596,-0.000492935172276221,0.00909197461221201,0.0129267549760068,0.00970825786285956,0.00936037441497661
"3446",-0.0173637191102232,-0.0135850794381763,0.000519283365068235,-0.0160561506997705,0.00508268208666229,0.00123285939398121,-0.0133934011044271,-0.0143979205802336,-0.00322314116542255,-0.0100463678516228
"3447",0.000509116017106237,0.0102707516339868,0.0129757787712073,0.00965299975421741,0.00213240108047263,0.00155969463142336,-0.00555340800933823,0,-0.0000548613373668738,0.00702576112412179
"3448",0.0131712565246371,0.00231058230847014,0.0071733903872484,0.0161620532665605,-0.0000607672680147386,-0.000901565430676765,0.0268055683495096,0.00830017572705133,0.00789258439943952,0.000775193798449703
"3449",0.0050523962414879,0.00691560611075137,0.00457861616790534,0.010528718873851,-0.0024320179824161,-0.000492255939421593,0.0116026480441818,0.0125122590799907,-0.00239274567617997,0.00542215336948115
"3450",-0.0039686553335907,-0.00114466575091576,0.00354488509301532,-0.00133012632830576,-0.00298656048695112,-0.000574515777232887,0.00537636424841637,0.00910578448927057,0.00283458167622652,0.0184899845916795
"3451",-0.00879520186967264,0.00229197794425895,0.00117744320979907,-0.00399556057703798,0.00305660834996191,0.0003284963536625,-0.0187760607673129,0.00515628776022314,-0.00548999290378871,0.0113464447806353
"3452",-0.0115127097360278,-0.00914699291104493,-0.004368313172043,-0.00780028989971671,-0.00310820937215739,-0.000903053951285648,-0.0215573960747999,-0.0182751044095527,0.00131170742685871,0.0044876589379208
"3453",-0.0111295722570011,-0.0309254543768542,-0.0148497642541264,-0.00920932165318966,0.00507420043088946,0.0018077321727461,-0.0278499606477897,-0.0254027873875655,-0.0200872983638749,-0.0245718540580789
"3454",0.0101843807988977,-0.00261969504073845,0.00308324763475087,-0.00748134192969074,-0.000790693459514324,0,0.0117137492086719,-0.00202839756592288,-0.00484631228060806,-0.00458015267175571
"3455",-0.0231909575485664,-0.0126552766796735,0.0058060279063179,-0.0155322296832395,0.00133926459270062,0,-0.0287538004550285,-0.0162601287262872,-0.0216064994662132,-0.0115030674846625
"3456",0.00266546293087666,-0.00169284167800932,-0.00390499137843836,-0.00464027863759986,0.00382995915162132,0.000492167002824173,0.00443232961064188,0.00550964168355228,0.00371879985143075,0.00465477114041879
"3457",0.0161669582689334,0.00145351263211047,0.00153400380207969,0.000932330958865579,0,0.000819798307432285,0.0202465663758638,0.00445202039547876,-0.00284997716769297,0
