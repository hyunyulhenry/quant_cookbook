"","SPY","IEV","EWJ","EEM","TLT","IEF","IYR","RWX","GLD","DBC"
"1",0.00212211723093758,-0.0056814470354658,0.0105634486272226,-0.0138089777070859,0.00606370035074288,0.00362855334275047,-0.00023823488591701,-0.00743695293540392,-0.01011555892928,-0.0260503050587256
"2",-0.00797621060863463,-0.0147621811294277,-0.0257840791300752,-0.0292382644144845,-0.00435303561055334,-0.00325411447288704,-0.0155038356414278,-0.0124338834144747,-0.0240065523436642,-0.0034512995305368
"3",0.00462525850329132,0.00164362834500564,0.00572253572691861,0.00725719012180659,0.00179375342128152,0.000725508719865431,-0.000242291002061856,-0.00339005251821212,0.00515210254785115,0.00519471605092869
"4",-0.00085063404212915,-0.00376383560049154,0.00640105341404884,-0.0223361655072509,0,-0.000242051126348675,0.0117532828011679,0.00161984607578791,0.00611769179894184,-0.00861317890472024
"5",0.00333218590726614,-0.00561872122315621,-0.0148410172356069,-0.00230329759424897,-0.00447655817073112,-0.00169152685184759,0.0159283875061749,-0.00565973401716846,-0.00427276924479103,-0.0147698688123383
"6",0.00438034628578832,0.0108136598205906,-0.00502142829521812,0.0126501433345514,-0.00584330071208583,-0.00266285792304721,0.011434232773009,0.00325225341279767,0.000660191450734482,-0.00132265790941177
"7",0.00759764933177887,0.00905914380438233,0.012977654262998,0.0203336969156163,-0.00463593496080827,-0.00206340397280125,0.00349644318156694,0.0066461799883657,0.0253999171136414,0.0233996224013486
"8",-0.00195494125685913,0,0.00355853205057222,0.00357477449165522,0.00215855100726814,0.00194603168953456,0.011498551045364,0.00257662121805935,-0.0032169375331168,-0.0228645994088241
"9",0.000419285258396185,-0.00057304824329707,0,-0.00418516439316152,-0.00306132541125947,-0.00194225200558251,0.00298488316759649,0.00706691963382089,0.0108116506243077,0.00883002834000157
"10",-0.00335593824303038,-0.00305809478065688,-0.000709148162663986,-0.0105519514238314,0.0030707259024958,0.00133804302799878,-0.00343395395127677,-0.00111633312218817,-0.00606642729991103,-0.0105032427762808
"11",0.00196434131967727,0.0107364911411358,0.00709716327695142,0.0179850132533814,-0.0027208412501557,-0.00157946327278835,0.00884491489780159,0.00974008347589694,0.0118856733660673,0.0150376039605462
"12",-0.00308061133924431,-0.00701852575518147,0,-0.00115424583911428,0.00238666131318577,0.00182497404382853,-0.00307406491442341,0.0102782122775675,-0.00444442857142857,0.000871366900456527
"13",0.00294968074128277,0.00897792590611513,0.00563793367584275,0.0227532330831659,-0.00657599298036859,-0.00291473823253452,0.00285569117551665,0.00751301689480566,0.0240752866059424,0.0317805604448693
"14",0.00805291846133138,0.00511179600558109,0.0133145799163663,0.00869061932587689,-0.00011381655425613,0.000122195086190935,0.0136673611919413,0.000931725508000136,0.00155688923134556,-0.00843882505047222
"15",-0.0117402782296068,-0.0154451339250472,-0.0165973490401511,-0.0307572789044992,-0.00719075986827777,-0.00389693993514073,0.00595544773789891,-0.00589752823026901,-0.00419717070737846,-0.00893599478055107
"16",-0.000913719080819275,0.00277388619729968,0.000702927752839422,0.00613326450503893,-0.000805198974248023,-0.000121490792450274,0.00301540518920729,-0.00624502224335111,0.00171714023469072,0.0124515654514379
"17",-0.000562421996066487,0.00228937836540988,0.00351375549550559,-0.0132524430965038,-0.00218642432945881,-0.000733995188640924,0.002894823826598,0.00612686175776944,-0.00623341144564171,-0.020356203459988
"18",0.0052092580776697,0.00532981302560187,0.00630267383024541,0.0154896664835846,0.00115304517504278,0.000978686116337002,0.00344275911189351,0.00405980399307748,0.00705662537243201,0.027705554222162
"19",0.00672302397912539,0.00511194143821414,-0.00417532450434566,0.00775909297911315,0.00840836710592052,0.00366662620902414,0.0113973055211385,0,0.00949861399099006,0.0105308029970261
"20",0.0059826595137642,0.00781788600721289,0.0132773618769466,0.0122480189860927,-0.00120482293762592,-0.000721164785794426,-0.000547169583573592,0.0113531482946263,0.00601571784619104,-0.00375161049023653
"21",0.001383086123111,-0.000934605986404935,-0.00620689907498195,-0.00302503939292709,0.00126349866742426,0.000856889977828956,0.0071156124208327,0.0110719997552913,-0.0144127872675132,0.0129706315284444
"22",0.000276393574802025,-0.00327423655290127,-0.00763353448627713,0.000953849250799887,0.00137627403694629,0.00110051350399898,-0.000651970773024146,0.00304159738051824,0.000466692602157481,-0.00330437818714768
"23",0.000276101252362437,0.00656976193527181,0.00839171797977034,0.00987340000263726,0.00549694060029648,0.00280724020913303,0.0137043244951343,0.0103107482538214,0.00746389387230284,-0.00497302215289619
"24",0.00220871307203674,0.00372976539313519,-0.000693643549549372,-0.00385930099273324,0.00296103493409827,0.00219199277163096,0.0146999253164435,0.00405259749277564,-0.00246957860056218,-0.0120781760068096
"25",-0.00130855480968306,-0.0023223791723983,-0.0124914998459981,-0.00533792453258242,0.000795520563912522,0.000243195786732153,-0.0076136368225258,-0.000597945128866462,0.0137706953630217,0.0231870629732278
"26",-0.00744727127439004,-0.00595931686280271,0.0028111715201582,-0.0119449851553155,-0.00567377314296436,-0.00303682085389001,-0.0141714245657776,0.000598302881159807,0.00915760115190478,0.00618051849681645
"27",-0.00340431820190334,-0.00327819738511537,-0.000700785356489764,-0.00683301014310367,-0.00228204481096439,-0.00134005522646685,-0.016753321842907,-0.00822091221572008,-0.00680588293379225,-0.0188371198035659
"28",0.00843510936031744,0.00977352256735409,0.0210378336471537,0.0158771923118854,-0.00217343798234815,-0.00073157249174105,0.0178078952457128,0.00813838248220544,0.00258867070469515,0.0183639546801622
"29",0.00656696595404482,0.012843145344263,0.016483502561536,0.0215332804796007,0.00951445412387897,0.00573773868404026,-0.00615606155632598,0.016594535325928,0.00804992454738307,-0.0135245569450847
"30",0.00130516637973477,-0.00202127542937802,0.00810796746504328,0.000594920337946947,0.0029518353564455,0.00157763754521612,0.00825911512155364,0.00294107174111069,0.00060269697441484,0
"31",-0.000480540638432947,-0.000276345719207538,-0.000670091816536211,0.00229403426731922,0.00350965175226192,0.00109104189329612,-0.00344888404107513,-0.000733162437638546,-0.000752943788408844,0.0174491644849777
"32",0.00212746561272059,0.00349958807310791,-0.00335342141618133,0.00262722434384988,0.00225588811972632,0.00121067659451723,0.00843618704890825,0.00190777150778976,-0.015822829779644,-0.0110249158425911
"33",-0.000411120809875043,-0.00734191770007731,0.000672961455531862,0.00295815791524867,-0.0016878310096945,-0.000121455803772319,-0.00525540417835391,0.00322172408437393,0.0312356463400902,0.0214698305811687
"34",-0.000753510666783752,0.00286603530410812,0.00268993301217724,-0.0025284473772873,-0.00541209558079148,-0.00253880231451831,-0.00506732252874265,0.00627747419464986,-0.00296950268654794,0.013742936552138
"35",-0.00390735909267936,0.0025814158309363,0.00871910017145616,-0.00718192335541168,0.00714143028365943,0.00400129527500748,-0.0141960601912247,0.0068182194260864,0.00848844352975586,0.00637963267720099
"36",-0.000894673435136384,0.00505723257650148,0.006648870663025,-0.00042540488468068,0.00664170669752928,0.00313954835913011,-0.00648532923077749,-0.00806879490540724,0.00561129643220171,0.00277337747782158
"37",-0.0390576856400801,-0.0539797589651595,-0.0237779997195946,-0.0813112101773937,0.0126352532668017,0.00842648023561199,-0.0324192133334843,-0.0368973165207505,-0.0395006472687415,-0.0189648488774585
"38",0.0102507808323093,0.0135396929246925,-0.00135329040260435,0.0250231500191431,-0.00452696626813109,-0.00346178051197665,0.0077761171697972,-0.00558084596516895,0.0163583387030521,0.0153039919303792
"39",-0.00298045563218152,-0.0131677865761087,-0.00474243921543993,-0.0143761011824965,-0.000634746113057472,0.00090078148277617,-0.00624080434063523,-0.0121339830995065,-0.00992784251228152,-0.00713994426755238
"40",-0.0130951163938767,-0.0130538223423906,-0.0163377949158395,-0.00926534596875328,0.00501347852285594,0.00324343096067992,-0.0206667998469435,-0.0188852219444052,-0.0320571406867212,-0.00918906513063011
"41",-0.00951868191508998,-0.0202802726485757,-0.0145329208160516,-0.0256479890148159,0.00166289542962317,0.000597467858420631,-0.0354436632604923,-0.0228483016595444,-0.0122429604809757,-0.0149191936410714
"42",0.0171095733899342,0.0276002791959264,0.0238765807448114,0.0439036793773289,-0.00298737802822169,-0.00131580931245812,0.0344495887428959,0.0281872961961696,0.0193866518353727,0.00941465989397505
"43",-0.00100205817221699,0.00194630887603853,-0.00205771841604041,-0.00609923213466057,0.0038845905160183,0.00179688328244887,-0.0142556740253735,0.011837646699947,0.00233828519600054,0.0137874316339257
"44",0.0084549776934546,0.0103921203866397,0.00893474676034223,0.0258288264705291,-0.000884824140326645,-0.000119561793025413,0.0160032402640675,0.00369463347045684,0.00279937778540984,0.00160000109706515
"45",0.000284164231645789,0.00288392299807483,0.000681296107118534,0.00178612247356358,-0.0105140257113004,-0.00562022627224079,0.01224984982925,0.0111963101287289,-0.00356704387870443,-0.0131789655455684
"46",0.00149177863631866,0.00383404043896163,0.00816876254923216,0.00490160926474981,0.00391486448805511,0.00276571062076569,0.0050715719648744,0.00712858898428381,0.00186775097276271,-0.00930789262729326
"47",-0.0194343898655909,-0.0244437308822566,-0.0182309316812997,-0.0290906946734778,0.00601693035751216,0.0044370833598355,-0.0263756097939822,-0.0191262290580164,-0.0100979022791097,-0.00776139923920816
"48",0.00745045644582132,0.00371937922979915,-0.00894089108085183,0.0082213996463949,-0.00454124721249571,-0.00131392832273791,0.00471106853105407,-0.019653034104846,0.00345257370601737,0.00205841743606472
"49",0.00136426859552419,0.00477789241622006,0.00069412502489552,0.00815439476960855,-0.000110856139938553,-0.00107517830461101,0.00750279529168463,0.0117463059024152,0.000625602136778314,-0.00616274323701982
"50",-0.00280017801508137,0.0034937961555106,-0.000693643549549372,-0.00853801249608155,-0.000223347783929295,-0.000118841942835846,-0.00558513266724336,-0.00346399722968183,0.0100031728665209,0.00248040983341546
"51",0.0120552510214507,0.0149904973330299,0.0111033767470741,0.0219365530068458,-0.00211396977525069,-0.00131811412702487,0.0100631171226238,0.0194856900498053,0.001856932751922,0.00494845688755019
"52",0.00549204406095005,0.00981403388292557,0.00892248211239877,0.00656378045720207,0.000557120736522254,0.0014388667855838,0.00324396594962439,0.0151375034270091,0.00818657733044725,0.00123089067396864
"53",0.0164579325687493,0.0245329850795801,0.0108843511171168,0.0299607704452685,0.00044626540558701,0.00143573148041809,0.0140870985853083,0.022744027385436,0.00842658227791837,0.00163947728165459
"54",-0.000768147492436366,-0.00653891912286053,0.00134584084009148,-0.00427785120718527,-0.00791096900943711,-0.00334551496976265,-0.000796550299791532,-0.00589075828087504,-0.000911546642357819,0.0163664913648924
"55",0.00146664528930995,0.00519146589935993,0.00134417541811938,0.00464005703573256,-0.00280849003008132,-0.00155921064037634,-0.000264161683275366,-0.000444534846241296,-0.00927615543564009,0.000402619932218462
"56",-0.00132510767416527,0.000737451822004243,-0.00536936136791577,-0.000598567991106691,0.00123887217096796,0.000840484205572922,-0.0155084745713523,-0.00340895554770126,0.0105908515551543,0.00442656260043939
"57",-0.00237437398209239,-0.00608222956638382,-0.00404840025328812,-0.00445030411881486,-0.00168585587766856,-0.000240352557684287,-0.00828457979881914,-0.00654354479643604,-0.00212635189102994,0.0028045321486756
"58",-0.007279582176833,-0.00917954572881796,-0.00745252251999162,-0.0178804558497069,-0.00202866592564777,-0.000119000273863024,-0.0116482854041269,-0.0074851487934916,0.00532733662073093,0.00958850037405323
"59",0.00105756347506825,0.0103874095163914,0.00136504946009786,0.0198690166944311,-0.00135451211461868,-0.00144124457602302,0.00535719258879697,0.00829582094660819,-0.00605603303303415,0.0193905524746216
"60",0.000211386171609984,0.00342710258784806,-0.00681656670538833,-0.000171371992107483,-0.00192277927212103,-0.00120183482071379,0.00935399353587885,0.0127149316368758,0.00137084535046927,-0.0147516879941152
"61",0.00112660002024079,0.00359983160951161,-0.00549089021858618,0.00686667714845512,0.00165970307821905,0.00111187490724296,0.0118495306774409,0.00531746809779121,0.00167325834113963,-0.00985019969883938
"62",0.0107627621057,0.0129679101795244,0.00828170462817934,0.0163682063322272,-0.00124780124190382,-0.00084443707943882,0.00869545927963444,0.0057302194227411,-0.000303659842176507,-0.00397922538928086
"63",0.00111376510255257,0.00254208637838649,0.00752926702828605,0.0062908471932468,0.00102162167007958,0.00156940990788068,-0.0065515847010531,-0.000876816792778179,0.0148867684980474,0.0111865837697289
"64",0.00271094059807253,0.00443776074955826,-0.00271750944657612,0.000917149464970235,-0.00374555180114489,-0.00253161334132546,0.000809371080963794,0.00438655120670339,0.000748435885299825,0.00197546276217331
"65",0.00138637569898514,-0.000991871460438332,-0.00136242605965198,0.00574623482636394,-0.00660972555704731,-0.00459553615926345,-0.000693508254165698,0.000145487216706597,-0.00493571634855339,-0.0102523310478511
"66",0.00117690067112575,0.00722028807430797,0.00341077438500492,0.00471954668250496,0.0029829359331599,0.00206546124743112,0.00254514789899529,0.00611381055625571,0.00946948759160504,0.0139442326305543
"67",-0.00407973881943935,-0.00394250357155157,-0.00407892131244625,-0.0092301576480246,-0.000686560521510393,-0.00121193712358347,-0.0133855633769285,-0.0111397069973358,-0.00119121493798613,-0.00157179448515576
"68",0.00444381578622277,0.00710665171022273,-0.00136502864824439,0.0167192972759918,0.000228426043272334,0.000970547485096285,-0.00526275532068343,0.0055595223456617,-0.00134174116452757,0.00590315003881492
"69",0.00456231264337204,0.00741413958928616,-0.00820251320691545,0.00490890979360059,-0.00308929697105886,-0.00169780058860414,0.0109350308863136,-0.0033463457397529,0.0126884314879365,0.00547739648670853
"70",0.00949615770434753,0.0117039976117963,0.0144728881349361,0.0118861717016479,0.00550958182031502,0.00109344884422824,-0.000233220243258558,0.0157662414411588,0.00825480591125038,-0.00778202330855171
"71",0.00265868251900003,0.00131475184029761,-0.00611404931401727,-0.00539078088836098,0.00559388041581332,0.00424567755055283,0.0143092620321452,-0.00546132976587088,-0.00584798228514671,-0.0101961268708496
"72",0.00122370079019252,-0.000525043946775883,0.00136689449839378,-0.00744194304197887,0.00499442957873053,0.00229510602382121,-0.00355599769166326,-0.00173388857020862,0.00558819117647058,0.000396154335922549
"73",-0.00027163739025593,0,-0.00477813097111568,-0.00806830304201334,-0.00169433770376759,-0.00012012726056998,-0.00863217710415964,-0.00376364425656672,-0.0124305065412623,-0.00277227922738532
"74",0.00944097433774815,0.00796903061946175,0.0041152068025827,0.0119132133174236,-0.00260255021632616,-0.00108470737721056,0.0109138345829609,0.00624801483188464,0.0173256036920717,0.0138999306258629
"75",-0.00376805638937483,-0.00564732072804763,-0.0109288753716594,-0.00397851200956556,0.00363086494968679,0.00205124693193715,0.00849890122609898,-0.00216667578191976,-0.00640458543251454,0.00665883749617335
"76",0.000405382914122843,0.000174717471578711,-0.00138139130624471,-0.000162971292866132,0.00372969871592521,0.00192677109069295,-0.00683340085736051,-0.00723569616177533,-0.0077644152427655,-0.0136186866940441
"77",0.00918170724853895,0.0105704404061056,0.00553257619194913,0.0123928979787151,-0.00349017845448463,-0.000600261088616327,0.00137638090962189,0.00918379599978092,0.00236226181770594,0.019723922310988
"78",0.00113694129234387,-0.00311165505497513,-0.00481430015824069,-0.00265772136689901,-0.00723331106737002,-0.00288723323685725,0.00137367909129993,-0.00548928169411622,-0.0150242453236743,-0.00696329557888986
"79",-0.000801423102020249,0.000259700014310527,-0.00552858371672771,-0.00500646041669217,-0.000226596528522083,0,-0.0033156262914501,-0.00072540296165946,0.0103184532532472,0.00506419748851039
"80",-0.00829292241092483,-0.0039009217342838,-0.00764446072803826,-0.0193147833762282,0.010474112343108,0.0043424688620004,-0.0191602244158691,-0.00218053254612749,-0.00695680896852591,-0.00891469419041446
"81",0.00256278364702744,0.000261036847139851,0,0.00397206159562646,0.000724022675197666,0.0000484715620463483,-0.00526366472232132,-0.0033504460081093,-0.0059620513317663,0.00195550177609105
"82",0.00585175024652451,0.00539449858300833,0.00560246451473922,0.0198646892151604,-0.000565390486116146,-0.00120569251388336,0.00823079612442457,0.020169738063972,-0.000449812552112516,-0.00780644828912236
"83",0.00541666555618492,-0.000865322462401452,0.00139270147481896,0.00840553494981022,-0.00226126714172048,-0.00108617933979149,0.00396568997043745,0.00286527365188971,0.0124511543683676,0.00472082218868608
"84",0.00379130584227383,0.012126497658171,0.00347718702147004,-0.00032058179557215,0.00407976357766771,0.00253803801324648,-0.00499532398856273,0.0062857662642779,0.0103719665245805,-0.00195784038455937
"85",0.000198721286754688,0,0.00485082990224139,0.00649425440611129,0.00270873483686507,0.000842887070641396,0.000933899875267485,0.0052528071153648,0.000879865057050289,-0.00470760579377849
"86",-0.00132534231480819,-0.00898608348890595,-0.00206892430402872,-0.0129840919289171,-0.00225159120859475,0,-0.00653208369238123,-0.0121455168147236,-0.00542128937728936,-0.00630683405612698
"87",0.00271984006788561,0.00276386397667649,0.0124395346054402,0.0161406542820308,-0.00394833633812586,-0.00325103262008852,0.0116241840311404,0.00114383194778744,-0.00633470858874685,-0.00515664530307158
"88",-0.0104522571962546,-0.0201518831413005,-0.0150169384552497,-0.0244616730670175,0.00237906732734094,0.00253652736300891,-0.00998166166425396,-0.0075679651217595,-0.0214973619643007,-0.00398732915969924
"89",0.0085575239707476,0.01687440920081,0.00762286853376204,0.0254005686869998,-0.00350354949147003,-0.00204826023844173,0.0111373936285142,0.0141005387400455,0.00681813636363637,0.0148119473263204
"90",-0.00218776707981516,-0.00216048906061439,-0.00275106760484156,-0.00992458799659701,-0.00260827690647447,-0.00144953437252304,-0.0104351916260709,-0.00397305479865939,-0.00255828453987728,-0.00355029840873888
"91",0.000266082325628414,0.00259834422849736,-0.00827582337901067,0.00120306029185691,-0.000341098233857529,-0.000120767709184122,-0.0134738177805481,0.00284903229767908,0.00392278219557607,0.00989703519012286
"92",0.00684058261710052,0.00216006846614691,0.0020861892376951,0.0144975472101769,-0.000681663119086795,-0.000603794344530395,-0.00926381447623847,-0.00724386632084262,-0.0141268858712521,-0.00980004381165411
"93",-0.00197893278444938,-0.00172436592431247,-0.00832759603573918,-0.0036321094714088,-0.00409701071530078,-0.00266313573273846,-0.0179812116278759,-0.00887131965103782,-0.00823170756803993,0.00831350277362031
"94",0.00872399814013325,0.0125218186465905,-0.00279919708628318,0.00515096712373531,-0.00662793110312765,-0.00291206569894742,-0.0086668727393131,-0.00389776103149653,0.00707038140394678,-0.00157051832110122
"95",-0.000524103143328514,-0.00759071203903516,0,0.00181347295366008,0.00299122137883079,0.00133912382781221,0.00689558414085956,-0.00130427117531928,0.00228939265671824,0.00983104263365253
"96",-0.000786639296942115,0.00120299786015798,0.00982478733076642,0.000157131367967578,-0.00516136252292421,-0.00279474056685314,0.0103955360683152,0.000580119218223318,-0.00715701255236845,-0.014408109306017
"97",0.000131267965503445,0.00472108868529797,0.00138971318578474,-0.00157380044134237,-0.00288224460934361,-0.00194994886194111,-0.0078680547936627,0.00203076588208373,0.00521478551601784,0.00474108523167938
"98",-0.00905262184544853,-0.0105935130299306,-0.00485764798255295,-0.0240348196359494,0.000925360244977913,0.00134292393027868,-0.015249144931332,-0.012302696186246,-0.0120537227333885,-0.00550522883832627
"99",0.00417049143404924,0.00682151114313778,-0.00418431437043032,0.0153415728567659,-0.00231076902858085,-0.00109693112705322,0.00631787948062601,0.000292604905226979,0.00293439382239402,0.0122577335130811
"100",0.00362585442305918,0.000428523135259873,0.0105045062029749,-0.00341990802406034,-0.000115971577586693,-0.00207519846302207,0.0305308629376244,-0.000585499557821723,0.00200181700025182,-0.0218748918446232
"101",0.00814458538086504,0.00488654191842497,0.00207879127072053,0.0102140010549032,0.00208448896556135,0.000978569869939383,0.0255642655142876,0.00630296731393964,-0.00537880743814345,0.00958467109811956
"102",-0.0010420115769928,0.00153572926680678,0.00968176585477165,0.00284362258960669,-0.0018487172811319,-0.000366628203002151,-0.00267893548519749,0.0180628643881442,0.012669962721416,0.00909802267606286
"103",0.00495676694062586,0.00894358011399699,0.00547960824917082,0.0249687085141439,-0.00525327962137223,-0.0043082011478579,-0.000466965996479884,0.00300431941432633,0.0137320870654245,0.00744810721222477
"104",0.000129845306391596,0.00303946401832511,0.00340587822522154,-0.00445687779336734,0.00455726071314988,0.00160229184731331,0.00630953466399564,0.00699002562223927,0.00150510230267598,0.00894950605841682
"105",-0.00395832290287146,-0.00547107483769249,-0.00135755316700314,-0.00347406071131062,-0.00628118305837932,-0.00320086503906458,-0.0173014798797931,-0.00878279420648764,-0.00255482412752006,-0.00385662185426483
"106",-0.0107500589535405,-0.019803797772653,-0.00407892131244625,-0.0251740576099074,-0.00046814782350435,0.000494094064061423,-0.00626223174540141,-0.0195802684858266,0.00060269697441484,-0.00038718847866448
"107",-0.0180453515461212,-0.0231391551176165,-0.00409543974624027,-0.0154153122701323,-0.0179152157440348,-0.00999576527446477,-0.0309157919837248,-0.0236148120264048,-0.0173166982492577,0.00503486046064849
"108",0.013011606842632,0.0142301890291019,0.0047976128104803,0.017674317317683,-0.00083510994138547,0.00186976429748298,0.0164415347049791,0.00104502662887573,-0.0159362698150086,-0.0177263688049796
"109",0.00172148171213515,0.000435819810067795,-0.00136418080851974,0.00856453686221914,-0.00286360883612213,-0.00261254123361665,-0.0147267374424296,-0.00372845905648733,0.00747424466717161,0.0192232805596453
"110",-0.0109059951354826,-0.0164634976537413,-0.0129782438596471,-0.0173769193330072,-0.0144815457851105,-0.00711084344785529,-0.0210732199493551,-0.0176644848560924,-0.00927355529861917,-0.00269446454548161
"111",0.0149687173985951,0.0172704617003778,0.00276803372271828,0.0200049487879173,0.0119013223510427,0.00326630886994606,0.0215268602093661,0.0118865774800763,0.00670828414066427,0.0127363633446651
"112",0.00638597500190974,0.00948964812643371,0.00138045945190224,0.0156895346495765,-0.00252038445727309,0.000250634339427735,-0.0102916949028838,0.00135522326459991,0.00108475129528518,0.00952748724430674
"113",0.005689991865653,0.0125055414391109,0.00895937692259241,0.0227855180651497,0.00685762950480662,0.00438217215085945,0.0151027635000887,0.00811302965534311,0.00386996916006099,0.00604001949708444
"114",-0.00117561913493547,0.00212927936610474,-0.00204928518371184,0.00090597809933346,-0.00203137471702675,-0.000498509898972488,-0.0148780636238386,-0.00330937739757875,0.00154200467361609,0
"115",0.00248519617560894,0.00144504543524793,-0.000684560398927059,0.00113201455145151,0.00933968789876416,0.00486321369281772,0.000990368731327296,0.00739490382359964,0.00816021592733862,-0.00975602421892541
"116",-0.013897423997743,-0.012985987630718,-0.00684916573980365,-0.00851659384496517,-0.00806744087792644,-0.00322605242849194,-0.0178083748234368,-0.0112359133623741,-0.011759376370218,0.00113671378480618
"117",0.00555765548642473,0.0061054674010339,0.00482756013323149,0.0124661661078524,-0.00478319473933098,-0.00124559852599049,-0.00402977750804101,0.00378784487194017,-0.00231804979629191,-0.00454197639049791
"118",-0.00940897718217515,-0.00965825249949781,-0.00960858704466394,-0.0132132299356579,0.00648894818759138,0.0029925324655633,-0.00379255542230628,-0.00981140398379865,0.00340769837074673,-0.00228145187285711
"119",-0.00478255599973276,-0.00276163075156577,-0.00554407726304174,-0.00760804924166769,0.00549168201801709,0.00323178649940625,-0.0227156028967853,-0.0213410607810485,-0.00540288677682743,-0.0038110602241177
"120",-0.0102782270758831,-0.00519260263987698,0.00139365074198361,-0.00873978827196031,0.000237606345881103,0.000248492953330182,-0.00142835866365765,0.00233639053727197,-0.0125717988514669,-0.0114765510385546
"121",0.0142286745026776,0.0091346154839278,0.00208772590429351,0.0142307172884031,0.000949261447263483,-0.000124377782474872,0.0217165001076782,0.00310777451290911,0.000785900672522821,-0.00154803023238326
"122",-0.000132520294667926,0.00206890135442728,-0.00208337638544531,0.000228593610482442,-0.000236175133543792,-0.000619302896515461,-0.0039062174275114,0.00898534602451617,0.00926659366315663,-0.00310073611494466
"123",0.00033222571086422,0.00593606613352371,0.00974250871296767,0.00350701921699881,0.0103195856840346,0.00520616070436208,-0.00128984070057392,-0.00230314919838359,0.000155539988934361,-0.00077756390523942
"124",0.00904085930801379,0.0116309102547412,0.0179185857439246,0.0202841044573383,0.00525669480694124,0.00152294033073863,0.0251869739982631,0.0110805584739539,0.011669519760519,0.00622568534584866
"125",0.00362356801144958,0.006086572153992,-0.00203116583233764,0.00796731172658705,-0.00609715020465251,-0.00296634709359567,-0.00466151173525686,0.000456354391289659,-0.0043063520904193,0.00116001076655725
"126",-0.00105080183078121,-0.0034452067399634,-0.00271359525328907,0.00443229934836298,-0.0112066759710133,-0.00558003124298745,0.0160756357508043,-0.00654188403316713,-0.00494284846904058,0.00926999570093279
"127",0.00525721699931947,0.00758880000932982,-0.00476171305520023,0.0171359987729978,-0.00405598668738938,-0.00236831051120634,-0.00211771421868712,0.0124042760648453,0.00838250569334065,0.00841948881502264
"128",0.000784745347418347,0.00343098009555143,0,0.00968909069923241,0.00359402500016448,0.00362404097407021,0.00374540696342951,-0.00862215378695141,0.00646548655273227,-0.0022770415146578
"129",-0.0142394405428757,-0.0146774173466412,0.0020503521677413,-0.0196935724158199,0.0169490473629723,0.00684851154078014,-0.0304725942854716,-0.0122062862555741,0.00351795672306299,0.00722704709078603
"130",0.00709013787998947,0.0131183803760544,-0.00341067039671283,0.00825466619980375,-0.0103293160787526,-0.00346293236591966,0,0.00447980499785783,-0.00259105315361896,0.00226594368689348
"131",0.0157902616667172,0.0167086179038469,0.00684479010469952,0.0219534257246066,-0.00343908091237777,-0.00285427263341365,0.0125721949066446,0.0083037204264067,0.00886300400785434,0.0026375300692274
"132",0.00297928451089535,-0.00246509932357197,0.00475866207782749,0.0124070368972877,0.00273775016693301,0.00223981905400272,0.00950163736791887,0.00732078823488846,0.000151499552476508,0.00150315505542631
"133",-0.000128645212731038,-0.0023063048085098,-0.00202995623270441,-0.0098040566504235,0.00961274751868912,0.00397410032971934,-0.00552166644773988,-0.00408840713138825,-0.0031803574614625,-0.017636035275769
"134",-0.000516892857209905,-0.00132118349987298,-0.0054237383571436,-0.000777680718001883,-0.00211591838981151,-0.00210310234253608,-0.00643614315204766,-0.00881709646030249,-0.00106350653296861,-0.00611145817995895
"135",-0.00180924618874101,-0.00727507946593542,-0.00477170061118615,-0.0122442719389997,0.00376929779487645,0.00359432846178476,-0.00546145301852996,-0.00153361497119775,0.0132319847908744,0.011529517868204
"136",0.00388419599074363,0.0044135382650714,0.00479457890628354,0.00995971854253641,-0.000235219452357494,-0.00012353062181869,0.00332004548140596,0.00153597055864196,0.00585408259438247,0.00341949609782533
"137",-0.010124500824525,-0.0092029340989308,-0.00408994002323293,-0.00688182371236534,0.00903934370660409,0.00494149620847595,-0.0160379907098316,0.000766822442151316,0.00850619285162812,-0.000378725846339356
"138",0.00306164423544275,0.00317971831607222,0.00616022970577257,0.0289329062825907,-0.0016288173749367,-0.000369338222139248,-0.0174648918478698,-0.00766237865070873,-0.00162771525221317,-0.00454541746867632
"139",-0.0173413134320314,-0.0212712345598042,-0.00340132731618448,-0.0342291772159689,0.0037289194715231,0.00270574502158638,-0.0256748193159861,-0.020077261525553,0,-0.00761027412690252
"140",0.00204931770644112,-0.00196052603185892,0.000682524730049039,0.00575114056106818,0.00197321779250403,0.00134834649661708,0.00135128551796648,0.00315185608756474,-0.00844818425302818,0.00881890096296867
"141",-0.023679223570638,-0.0379159863285692,-0.0177352448100691,-0.0509649046240505,0.00834199453152684,0.00796043074934794,-0.0229419798200036,-0.0416341036443426,-0.0186846033278145,-0.0106421866674594
"142",-0.0196594551869486,-0.015178338242352,-0.00972227491988931,-0.012954847405439,0.00287173256168471,0.00194337704458425,-0.0276243251778049,-0.018688584845594,-0.00365571961444877,0.00960418518193684
"143",0.0156434395449339,0.0208198641982129,0.0168302797463482,0.0327355927746129,-0.00286350932870483,-0.00254615952440662,0.0134945506353523,0.00818573623780061,0.00550363825080957,-0.0114154519572044
"144",-0.011263316355819,0.00573948648774314,-0.004827412943186,-0.020466846675945,0.00723974410548611,0.00413325554875565,-0.0133148724153404,0.0122617719503222,0.000304150842518558,0.00808306373567436
"145",0.00487217797855521,-0.000527132112596362,-0.00762318547098906,-0.00392212131784686,-0.002165240649323,-0.00277120754911908,0.0156253302684735,-0.00965746132501188,0.002127967743913,-0.00152730162096215
"146",0.00798986503992638,0.00368897704491089,-0.00488834823728235,0.0110559869759697,0.00252481686229999,0.000730942594290518,0.0146850041436155,0.00495836133781813,-0.00060671924768696,0.0015296378393137
"147",-0.0257451141498606,-0.0175022068901207,-0.0140349519857694,-0.0431427138823994,0.00664069428638747,0.00645500235703289,-0.0368020086590932,-0.0149668287550782,0.0121414935823569,-0.0110728958450327
"148",0.0167596658551687,0.0115792673467332,0.0149465811135809,0.017847181292771,-0.0072786782271298,-0.00399255842337598,0.0260442065002695,0.00100141460274239,-0.00254918270957627,-0.0138994995789665
"149",0.0106693644396483,0.00255351676402493,-0.00210398007030288,0.00746009474834608,-0.000802329474432262,-0.00012217540806736,0.00404478589908019,0.0158469990154306,-0.000601232739081525,0.00548151681725861
"150",0.0139405114871491,0.0209028414607042,0.00843317174251856,0.0335876178754384,-0.0121538586007245,-0.0069260021701163,0.0362553113154673,0.0279146587674619,0.00436212375020517,-0.00155763343848836
"151",-0.0296334583001459,-0.0351858314956044,-0.0160280140095544,-0.0413586703520218,0.0013934353411329,0.00562828386691239,-0.00174296041184152,-0.0190096173578963,-0.0196195605640062,-0.00780031722738583
"152",-0.00467695404634783,-0.0141774257510432,-0.0141643410606317,-0.0173346848678908,-0.00231764004244306,-0.00145994441699504,-0.033167527728577,-0.00749088923157804,0.0169569357921926,0.00353769611988386
"153",0.00359326896837575,-0.00018105272980895,0.00143681150591668,0.00987884217664403,0.00290424838030945,0.00158354537746686,-0.00416695030368885,-0.0045940854917168,-0.00465672224725844,-0.00705053381947773
"154",-0.0152862310029342,-0.00986059503186076,-0.00286932510624893,-0.0258521117636407,0.00266356229672771,0.00365004224723031,-0.0376564299610854,-0.0214270644415084,0.000452746741540944,0.0031557362828909
"155",-0.0137749842789312,-0.0244859612151852,-0.0165468193363462,-0.0392895442146558,-0.00358028421452539,0.00181866572404532,-0.0108699885808752,-0.0296446834310861,-0.00241369735384378,0.00747162273480795
"156",0.0075154949808578,-0.00290345849685891,0.00219454294321286,-0.0170048850285119,0.0103182550931775,0.00387215482795433,0.0257877230082453,-0.0218713004883418,-0.0219264640220684,-0.0171741360556121
"157",0.0183674304791186,0.0186921664566109,-0.00729928810442637,0.0316451724158264,-0.00401673685353388,0.000722458076129362,0.0262823632507423,0.0216504079383144,0.00510207173778587,-0.000794281750049253
"158",-0.000484144058761848,-0.00138272763484171,-0.0110294840483774,0.00204524165095177,0.000576606222379095,0.00216767056493161,0.0167011762161171,0.000521308766866735,0.00169206270751987,0.00278215339106791
"159",0.00200519321744896,-0.00277043551796652,0.0126393287714133,-0.00367351937541505,0.00483524181371875,0.00432691702486565,0.0150583127703472,0.0111111476046293,-0.000767859301235019,-0.0015852880109033
"160",0.0118677860034349,0.0247224519941809,0.0132162028047402,0.0430152974192184,-0.00160388984237803,-0.0032313456911387,0.00809158029783963,0.0317648583112873,0.00507149223912728,0.00238181403621773
"161",-0.000886136310034868,-0.000813364266582739,0.00724630508698665,0.00510574975833911,0.00344298370611695,0.000360709421351579,-0.00709014933756491,0.00931928136165472,-0.00137620790898463,0.00316823425738266
"162",0.0123531180875305,0.0215227529857969,0.00503587786601112,0.0238376439223793,0.00492002430087135,0.000359496289690453,-0.0063325589862816,0.018961046336315,0.0122493190093194,0.0118436731577627
"163",-0.0093036255893334,-0.00894099627215661,-0.0078739609280396,0.00457994684368623,0.00523562669743161,0.00275890978845794,-0.0135592019561602,-0.00728137668399831,-0.0019663893213373,0.00117050424605614
"164",-0.021980428321395,-0.0241178535339428,-0.00937946155824454,-0.0406535234598203,0.00169883864018705,0.00514466890629017,-0.0316153363457701,-0.022167499821418,-0.00591098790947309,-0.0105221384053501
"165",0.0196214405994692,0.0259037942439122,0.00946826882168073,0.0396041688878754,-0.00271357211590384,-0.00380820373924184,0.0262597679709888,0.0218367814101683,0.00731825017949372,0.00945246275909684
"166",-0.00266112797279483,-0.0056212086793016,-0.00649368490666191,-0.00510437949228726,0.00668858821536467,0.00501672721640722,0.00484071582067314,-0.00897201448617868,-0.00408652943847421,0.00195096581230558
"167",0.00985279543412521,0.0171378171298595,0.0217863715832862,0.0258074331767095,0.000787781038423807,0.000238378181750765,0.0199587813815951,0.0139915814929996,0.0109421575558286,0.000389366640277888
"168",0.0100960469197986,0.00961550797941313,-0.00568552075851847,0.0168718028827097,0.00047419774278934,-0.00186083744901155,0.0134952279505887,0.0159088368274234,0.0138305027283752,0.0112884887874316
"169",-0.00865363907411387,-0.0139800689300233,-0.0192995932666494,-0.0151236413858125,0.00801727202555003,0.00621598364578868,-0.0239678772960406,-0.0209330920254038,0.0017793000658568,0.00192459985923144
"170",0.00230084314335866,0.00221555140549534,0.000728966992237678,0.00782713858132955,-0.00257685703371813,-0.00213828612793088,0.00613927577971007,-0.0052228342097741,0.01924220009598,-0.00384172346283407
"171",-0.0139068985450549,-0.0115826532923822,-0.00509856336470405,-0.0225592801875587,0.0141512293568633,0.0107145355646454,-0.0187122660093051,-0.0164070961965407,0.00769674691117128,0.00655603403984628
"172",-0.00191669621327384,-0.00581455922404506,-0.00878455482549201,0.000756844524342215,0.00775272890299927,0.00223870542787319,-0.0189304150015427,-0.0145117272542488,0.00331465633830019,0.00689651548866221
"173",0.0116605951357276,0.0197050166967021,0.0103398803051493,0.0201886583147695,-0.000769350752755305,-0.00211560806406341,0.0180284964510367,0.0189570294655603,0.0129272329965284,0.00228314746503155
"174",0.00257665994760869,0.0032648055133746,-0.00292419264096055,0.00355800918959215,-0.00373917265983548,-0.0024729529395201,0.00179837397856097,0.0101330902564032,-0.000850794137158162,0.0106301868737808
"175",0.00703302861264321,0.00562862121543861,-0.00733130684847505,0.011078410404276,-0.00894235734601556,-0.00590405881507949,0.0183680175034475,0.00970224767930739,-0.00539308835357777,-0.0075131534517725
"176",-0.0000678128790928545,-0.0099702948920718,0.00295424829890067,0.00197197858720921,0.00144857256356645,0.00130635776037957,0.00474582266683798,-0.00716589110164323,-0.00128430361631549,0.000757043374380428
"177",-0.00537223461472125,-0.0167841200482918,-0.00515463327301546,-0.00634234964657454,0.00478291556857657,0.000592618888842988,-0.00188929043553365,-0.0247705542045696,0.0140020435491368,0.0117245866427997
"178",0.0294395677546524,0.0420485978836016,0.0103626823733904,0.0484226914795836,-0.00752793642926564,-0.00106662799919488,0.0311023150709724,0.027754588280783,0.0102859798466115,0.00373824050057459
"179",0.00590320905270292,0.00353470064488226,0.0109890590984605,0.00454836983919282,-0.00925644477586374,-0.00356023062252242,0.0203275178230464,0.0193122342929073,-0.00376564869312324,0.0085661949880711
"180",-0.00704228219065572,0.0022338766914447,-0.00362306416853042,-0.0031347311915243,-0.0189126476374565,-0.0113155430650852,-0.0122106850173237,-0.00851001118655448,0.0180596528069437,0.0155096524025742
"181",0.00269857093620196,0.00642977559066926,0.00218150805111983,0.0132776673016606,0.00849084548593604,0.00505971598324284,0.000260013120915836,0.0131570702185018,-0.00522559123727184,0.00690905679580123
"182",-0.00184223681054174,-0.00170349933992853,0.00362850028397355,0.0124139087060813,0.00284514490405541,0.00131852010994171,0.00858610204188093,-0.00145190768555581,-0.000829375218654893,-0.00180574604944927
"183",-0.00197841983955394,-0.00392524837151398,0.00578460217340471,-0.00374675109116029,-0.00351766357960737,0.000119719485002445,-0.0165533708985753,0.00226194922373102,0.000691795803704931,-0.0072358181019565
"184",0.00528466683743312,0.00436890398461842,0.00862667071467205,0.0133335159140298,0.000910976252957107,0.000359066556065546,0.00569016067576711,0.0169243858553767,-0.00456244975632647,0.00145768792851686
"185",0.00591381811143332,0.0119402320091639,0.0228085047827999,0.0148446097940229,0.00693880951514858,0.00322952648093411,0.00947349784561302,0.0112534957641299,0.0097221805555554,0.0262008927706412
"186",-0.00333156306132665,0.00463553919553861,-0.00069687848834965,-0.00631665379914459,0.00225906399903342,0.000359390325865405,-0.00325854759107902,0.00705376962128423,0.011141747364859,-0.00319145367419116
"187",0.0112731230558929,0.0100670261063789,0.0111575125399204,0.03144861105368,0.00571487408667215,0.00119597854123454,0.0265464290613948,0.00498049765274033,0.00530540048142014,-0.0103167347210077
"188",-0.00136136583891244,-0.00299013800754522,-0.00275865685635202,0.00681179384911523,0.00315028075907375,0.00215153267672274,0.0091719420830525,-0.00263260849083657,-0.020974343140072,-0.0201293040553866
"189",-0.00201149422408331,-0.0036653071966819,0.000691640551272243,-0.0302837427053154,-0.00291667870575774,-0.000715459821345243,-0.000252458875563688,0.001552232481983,-0.00621970991623244,0.00110047505025279
"190",0.00156083888868053,0.00526756923347849,-0.000691162515249144,0.00996699379926258,0.00382530589031216,0.00178938763844405,0.000378679558013628,-0.00465079865904994,0.0134909731991384,0.013924485602435
"191",0.011881282085662,0.00756869085074019,0.0131397788432843,0.0333551752787224,-0.0107578448300295,-0.00881532014865638,0.0198157311837357,0.00934572153104307,0.0072732122708985,0.0028913363212475
"192",-0.00532538309638819,-0.011474390079083,-0.00546082219599131,-0.0106321697025316,-0.000792948030228002,0.00360589984811943,-0.0111383150437493,-0.0092591877408138,-0.0118529015843896,-0.0209009532259744
"193",0.00941746280493572,0.0125262560312283,-0.00274531955252999,0.0155725477185169,-0.00124701199959498,-0.00311328354246521,0.00575692856092802,0.0171338328406039,0.00772090180230101,0.00699301195640767
"194",-0.00166105613305678,0.00041245630274056,-0.00206471551512133,0.00133068296675587,0.000567467736789951,0.000960491141287712,-0.00136907298286515,-0.00137819332379718,0.00369414440794325,0.0116958755188288
"195",-0.00480089359430191,0.00412195715604646,0.00137948613179595,-0.0087954902821622,-0.00102088926338928,0.000120275987544938,-0.00672865678843748,-0.00398754802514034,0.00749731451066915,0.0111994302013048
"196",0.00553134043801906,0.00615771295669698,0,0.0182581608344197,-0.00488259252614354,-0.00335986431178159,-0.00727638406931808,0.000770347921683401,0.00920027010146018,0.00464463410506832
"197",-0.0084434061418619,-0.00873119834018177,-0.0117080616789698,-0.0122254824857729,0.000228067063543058,0.000962933679010902,-0.0205991342529729,-0.00846189339915293,0.00737368319472775,0.0170696735864164
"198",-0.00793496097767055,-0.0113599583306038,-0.0181186282276603,-0.0185340207238018,0.000342684111233948,0.0027663036352592,-0.0166452461382351,-0.0217219930903525,-0.000266116585921239,0.00104887679717081
"199",0.00305600456650512,0.0122396197606995,0.0014196274065017,0.0230872795735688,0.0109482394779432,0.006118419864928,-0.00275525544647626,0.00475821419739808,-0.00825350073535003,-0.00523930066369616
"200",-0.0036301469726524,-0.000493161428931188,0.00425211008107773,0.00505718235900465,0.00552809269209908,0.00381563099119853,0.00263157310772066,-0.00552511855827242,0.0201342281879195,0.0179073168434274
"201",-0.0261566758186695,-0.0198337524712986,-0.019759994230043,-0.0427675581404313,0.0149224298080344,0.00855223016107187,-0.0322832130186878,-0.0273014438426086,-0.00394740789473691,-0.00275953735000611
"202",0.00581284108846547,-0.00503802543375953,0.00575952700521576,0.00722743274676785,0.000109825062371227,-0.00188423965797335,0.0123401202163369,-0.000489681649533336,-0.0145310309589576,-0.00276717346854638
"203",0.00810427459412422,0.0156116832526456,0.00286331605762569,0.0277236218169916,-0.00132728029181439,-0.000236012617740422,0.00870754406414642,0.0179594047869576,0.00844510746501625,-0.00693725997684724
"204",-0.00184511640915996,-0.00124617849323672,-0.00428287454962073,-0.00653767605790867,0.00741667258730394,0.00507412385496453,-0.00398432951305783,-0.000160550005887439,0.00385476523243011,0.00349284216203993
"205",0.00237693863088051,0.00582366948441537,-0.00358395473917084,0.0127139193431693,-0.00340592001118067,-0.000821637655483487,-0.0026668158714962,0.013153698833789,0.0067532047174208,0.0233204754837524
"206",0.0117223849405106,0.0168733686694333,0.0172661709227624,0.0283262004676803,-0.00231453555612771,-0.00246829545503291,0.0147062431776979,0.0186825753325823,0.0218335265268121,0.0153063169226604
"207",0.00332012769819845,0.00618192787911753,0.0134369908488996,0.0230064055465338,0.00386683283018274,0.000824300071956774,-0.00724658470878325,0.00326429734363498,0.00553483059506155,0.0164152409450689
"208",-0.00694242985746152,-0.00727582582120334,-0.0048848306186946,-0.0188906239391676,-0.000550662332180818,0.00106010075110374,0.00451244953496155,-0.00325367637648222,-0.00985669444994774,-0.0224126033472398
"209",0.0103879436813026,0.0146580370246554,0.00701270386690056,0.0219437450420219,-0.00903006008615825,-0.00670226050597056,0.0179678632776168,0.0219148634152826,0.016418940308182,0.0283210275855652
"210",-0.0234073359334329,-0.0244780525440389,-0.0125349077734968,-0.0403734296779785,0.0129920630224627,0.00816169928439714,-0.0356910033762647,-0.0267677560949686,-0.00877643059871147,-0.0127869289061899
"211",0.00112536696707255,0.00822698204061978,-0.00282082543272433,0.00567216104827173,0.00319632950091586,0.00271008380028359,-0.0197845642163448,-0.00781354850127192,0.0243808802771717,0.0215875633978628
"212",-0.00760552034617623,-0.0134639589602653,-0.0169731102992449,-0.0347693525705844,-0.000439631094513615,-0.00117550648763731,-0.0142794542377161,-0.019530856688066,-0.00100215455337194,-0.00650202454672566
"213",0.0134620632714495,0.014061189658737,0.0115107879267731,0.0379477957054286,-0.0048353869529334,-0.00176503259708272,0.0104468866898546,0.00883499788667974,0.0210658307210032,0.0261779946862162
"214",-0.0273558045679061,-0.0160685751616176,-0.0184921031570132,-0.0318586007506626,0.00176752327519791,0.00365442711523944,-0.0337749341537441,-0.0195858127077254,0.00994716934790607,-0.00510201048791581
"215",-0.00507082079226051,0.00887016921766315,-0.0159420700350371,0.00511174065717657,-0.00176440464891403,0.00223149133266398,0.00627795738411341,-0.00357320618891199,-0.000121534536029588,-0.00256400139839019
"216",-0.0137261005499802,-0.0230074636117131,-0.0132550599377554,-0.0235220793747982,0.00850282883769626,0.00597564968190456,-0.00340305337090629,-0.0203750522339103,-0.000608087050659512,-0.0003214058130524
"217",-0.0099219243906471,-0.0159797958228595,0.000746193248328808,-0.055338617748541,0.00361351272036847,0.00174799711649865,0.000142760289126187,-0.0257898617221685,-0.047213397420297,-0.0218579729895122
"218",0.0304800342880163,0.0286323042383279,0.0171516258180291,0.070640893701329,-0.00370949919273544,-0.00511615987831771,0.0358462982089116,0.0401364195061542,0.0104725411057773,-0.0190600112852922
"219",-0.00276830708283449,-0.002907922456026,0.0029327686213807,0.00096552479408718,0.00109498786031037,0.00069995923265731,-0.0146938149947777,-0.0106737177237044,0.0146612229021277,0.0224454312693505
"220",-0.0144244696966345,-0.0166668674288888,-0.00877206530936858,-0.0230222564211353,0.00940758664822061,0.00560692292523446,-0.00557494661521507,-0.0182566579572576,-0.0290234433112039,-0.00982962716745794
"221",0.00171779583196363,0.00423735890730281,-0.00737489607814812,0.0123747487973558,0.0014087066681312,0,-0.0190608605473404,-0.00422658008158483,-0.00256570888642882,0.00330906930670882
"222",-0.0139241646366903,-0.0270040373328425,-0.017087458515992,-0.0460988745753405,0.00649239933106394,0.00720096509363088,-0.0191456735383004,-0.0280138049918582,-0.00655951125401932,0.00758579294261863
"223",0.00612104772962652,0.0222893732384184,0.0264551136382229,0.0274694643217368,-0.00107502904845835,-0.002652612210848,-0.0233064318109208,0.0155459905116631,0.0288710908563203,0.0248772327886559
"224",-0.0204641009867569,-0.0184947107678094,-0.0176733683470071,-0.0503518073806842,0.00581186989909432,0.00786200936490045,-0.0074572885223968,-0.0223596030413535,-0.00138417010967451,0.00127765068033292
"225",0.0172920456943946,0.0215228047988809,0.0224889755431115,0.0295495104461703,0.00299700677789416,-0.00298244380385171,0.0190834935264252,0.0362419474399132,0.0238155112926473,0.00925023354463761
"226",-0.022063266717857,-0.0197156590077066,0,-0.0396933255160701,0.0197375903357992,0.0136923569253842,-0.0376000558389396,-0.0290321511685323,0.000615421538461502,-0.0123260774232595
"227",0.0114935368342592,0.0125163116857656,0.0161290762428195,0.038295627060162,-0.0095217384470111,-0.00930721675365331,0.00735432307673478,0.0307742484244422,-0.014760208557434,-0.00800003976861519
"228",0.0319841211838172,0.032395627971058,0.00937954955064146,0.0547809002287301,-0.00675972515755374,-0.00355254055196497,0.0468442521640968,0.0154368363480824,-0.00661670428506134,-0.0122580734124823
"229",0.000339701274137294,-0.00908339034742622,0.00357412063628049,-0.0122583817324197,0.00861408830908506,0.00563387175432761,0.00799073833922592,0.00133660076617748,-0.016212152821415,0.00228622915887211
"230",0.0100560927333098,0.00374993324759165,0.00213627480086309,0.00849140201305798,-0.00485028934137699,0.00137280150147756,0.00922413002558731,0.00600596563290434,-0.0122636562629492,-0.0123820652419223
"231",-0.00659241863203164,-0.00356973706323627,0.00142166731415938,-0.00867886485765412,0.00793592405248367,0.0039529097620119,-0.00728304048013773,0.00364830224103674,0.0124159208484222,0.00725844226775885
"232",-0.00893841947936169,-0.00599911014930588,-0.0106458314714766,-0.00261346672342477,-0.000105498486802635,0.000912254814217306,-0.0261835986292704,-0.0133837977438539,0.0143076522011707,0.00458558632946859
"233",0.0167398537379027,0.00813033636826654,0.0186514443211649,0.0444125040982775,-0.0119282103156539,-0.00376248311439886,0.0285123830174574,0.0217719101230507,-0.00969779572549634,-0.00749915544072055
"234",0.0143136432094775,0.0106432339443117,0.0126760610556844,0.0157425812077283,-0.00875890951727343,-0.00526403181445723,0.0359094187889204,0.0136040439539389,0.00941124288736761,0.0180682734706157
"235",-0.000198595786302103,-0.00255058005367281,-0.0090404572675431,-0.0118554288381991,-0.0112081650449872,-0.00644249114701878,-0.00485308607877877,0.00258742335002871,-0.00970146114269388,-0.00322681525340973
"236",0.00775268204880875,0.0112174403718421,0.0028070545852994,0.0003123725231029,-0.00599456906683171,-0.00231556516587494,0.0250798996437254,0.00403241931475606,0.0178117307331229,-0.000647459196076228
"237",-0.027419580694604,-0.0268354472793245,-0.0216934520423043,-0.0423538026959146,0.0196266966718845,0.0136948472654037,-0.0572242276392579,-0.0224903216453195,-0.01450005,0.00874629264896143
"238",0.00987081973458026,0.0233846377821265,0.00786832850726782,0.0300065800351814,-0.0103233828314669,-0.0083575893642357,0.0031719190620465,0,0.0209284891389392,0.0272961382131933
"239",-0.00207558088673043,-0.0197377474614493,-0.0205817735031592,-0.0274857963272479,-0.0108662922645145,-0.00738982153104617,-0.0172468185533402,-0.0164334981089073,-0.0247235439116299,-0.0106282956909713
"240",-0.0126794349080525,-0.0252319824711406,-0.0391302905008757,-0.0238343651268929,-0.00461329103195951,-0.00290696029348381,-0.0302717532178629,-0.0342521960387819,0.000254738853503245,-0.00695106564738879
"241",-0.0142690026497956,-0.0173996515001944,-0.0173456162983323,-0.0426284500170245,0.00893854868866883,0.00594865780629439,-0.0180970550535446,-0.0501730914784668,-0.0049668876069876,-0.00489079563714301
"242",0.00558349614809428,0.0109911334849944,0.017651797606592,0.0274541672722677,0.00645426244540048,0.00197119143554625,0.0129011647727812,0.00273230699047056,0.0143351215026926,-0.00425944207669848
"243",0,-0.0101812337251252,-0.00678758402537016,0.00651120818455642,0.0132594031589219,0.00798630133631684,0.00833989374822997,0.00999024733820297,-0.000126208201892797,0.00954259968372395
"244",0.00630654174363254,0.00392273149096334,0.00379656263773898,0.00545770162214598,-0.00214504212008482,-0.00160726587047377,0.00375953403031337,-0.00629473879581544,-0.00719333688019519,-0.00423733058600284
"245",0.014415615812746,0.0145870394909495,0.0151284440555808,0.0301568659019555,-0.014619247272286,-0.00724592092914889,0.0170786725926964,0.0130326400469982,0.0181771963436428,0.0117839818799261
"246",0.00742548559909517,0.00679760470341573,-0.0016561270464257,0.0169132388094759,-0.00469012571657124,-0.00289648526460506,0.0272500694649107,0.0189190795170902,0.000499388277138246,0.00744093606279606
"247",0.00214447822155917,0.00550257946184884,0.00452475929424789,0.00518333649456926,-0.00876818032502069,-0.00476357507726588,-0.0166333188672757,0.01503032095503,0.0172198404943829,0.011881835103565
"248",-0.0125709723781873,-0.00277981780909575,-0.0157657196913448,-0.0230757794527133,0.0109014269937948,0.00671414098195156,-0.0194547830197084,-0.0243895941292711,0.000490689419431423,0.0034910490379898
"249",-0.0025057282311941,0.0083624485930256,0.0114417287112698,0.00376082974259884,0.0155938875384649,0.00803145193592036,-0.0147411610581255,0.0157140472572885,0.0176557385398661,-0.00316255885803629
"250",-0.00739978029586363,-0.0122668470739286,0.00226229999748773,-0.0120290131569113,0.00605621767573927,0.00461767672030544,0.00305356892231479,0.00123088039582764,-0.00650603614457834,0.00126896397825904
"251",-0.00875465259025587,-0.00271119474158721,-0.00451475038780724,-0.0165006262338848,0.0144022852922492,0.00712570320576633,-0.0083717508182416,-0.00438996741349196,0.0291050452231998,0.0275666024282257
"252",-0.000482957571239173,0.00175388613183647,0.0037795525084825,0.00899752046815827,-0.00137850382908622,0.0020542292117911,-0.0323866961032253,-0.00370365388520177,0.00836670977649412,0.00770883958221713
"253",-0.0245066454500248,-0.0234611337288972,-0.0256027168065389,-0.0300367093628903,0.000212774951478201,0.00261901295478095,-0.0317255454176857,-0.0219506561570099,-0.00514202407385755,-0.00581387407030654
"254",-0.000849092819244834,0.00502004387097243,-0.00618240969955097,0.00732701731362817,0.0043492086400243,0.00181683596959714,0.00933787655742857,-0.0162896976579424,-0.00422882664967084,-0.0181595601336975
"255",-0.0161481321164352,-0.0090983756862919,-0.00233257387666974,-0.00775398419664874,-0.00116280287679782,0.00215467708091621,-0.0363577633008321,-0.0220790850806291,0.0237112430238733,0.00909093024415042
"256",0.0105100383398615,0.00414108391558377,0.0218238322022217,0.032780035162097,0.00190418765830924,-0.00158387148120154,0.0197072369098492,0.00564447545392088,-0.00265033420892291,-0.00994093566611409
"257",0.00655413972607244,0.00080654537714353,-0.00839049364031019,0.0117850873317003,-0.0135092822013503,-0.00271902003538194,0.0132143855571809,0.00187044142195281,0.0196417901915036,-0.00470664262171938
"258",-0.00806842853002543,-0.0173774248952824,-0.016923188341543,-0.0281268698933901,0.0078100122753828,0.00636286763401772,-0.00163000887700371,-0.025209864515197,0.0037393994334276,0.00914241888765055
"259",0.00806271574164197,0.0165908766911871,0.0125194310083654,0.0147085456828111,0.00371528625883988,0.00045119897691448,-0.002776430743055,0.0153256382889604,0.0108376493376012,0.0124962089895626
"260",-0.0220128727210321,-0.0312948853451521,-0.0278207503687156,-0.0452318519054824,0.0112116486091516,0.00654532925163354,-0.0260355527526318,-0.0309432978279265,-0.0173107324401304,-0.0123419810154484
"261",-0.00861282931157614,-0.0216602871597643,-0.0182827229913249,-0.0416109231734758,-0.00721685660790228,-0.00190574967569201,0.012945433659606,0.00272600654945987,-0.0146607686023587,-0.00937191995711351
"262",-0.0259160811923892,-0.0142874774960327,-0.0137652874200634,-0.0291160514565815,0.0129582290321042,0.00808785995631611,-0.0121160887945434,-0.010874233724063,-0.002306770552714,-0.0129297788189532
"263",-0.0102675459089789,0.00105619261927825,0.0262725761660576,0.0228130963657633,-0.0068644505861809,-0.00144852844711751,-0.00840060236050311,0.0070674424750381,0.0106358150289019,0.00383388391305206
"264",-0.0101467217905142,-0.0312591271691831,-0.0368001830828457,-0.0251110742622984,0.0106816029725723,0.0111593448949565,0.0337174182732105,-0.0183235534974003,0.00857927267397107,-0.00350091581404965
"265",0.0240205967414078,-0.00653265262722247,0.00332235039548401,0.00636346992283299,-0.002279660771623,-0.00463521211144946,0.0817898008339717,0.012708539277676,-0.00317567206931324,-0.0188438187034397
"266",0.00844179833533065,0.0297896072831794,0.0165562700501978,0.019421961299356,-0.0200428266414496,-0.00909233021202815,-0.0195455669068106,0.028431545903852,0.0249175449416035,0.0247395512072714
"267",-0.0144454815795699,-0.0201239640770395,0.0154723926063782,-0.015211690906119,0.0168496223971646,0.00928832312600902,-0.0139078814628966,0.0285987014081639,0.00244228458165452,0.0222363674138357
"268",0.0165363928741649,0.0156991348390574,-0.00561323851586082,0.0247448081112029,-0.00375196646720577,-0.0036594483515624,0.0371413893875434,-0.00185371009656277,0.0160575520689628,0.00466139951663203
"269",0.00495406632347528,0.00767967676365577,0.0169351638415072,-0.00490249583913993,-0.00679983200247314,-0.00400471267468483,-0.00604431192944255,0.00185715271930942,-0.00653948773841961,0.0083512203980638
"270",-0.00735779604436926,-0.00347268800631062,-0.00475801954107113,-0.0131627287772461,-0.00653018495608915,-0.00044794562380257,-0.0234111804207492,-0.0157557721585736,0.00998349950667032,-0.00858889055647272
"271",0.0182341335873208,0.00948668547636156,0.0135459459602427,0.0200448985139179,0.00710354407558911,0.00514162451790612,0.0238169077317343,0.0169492675338891,-0.00716919415966089,0.0049505395663092
"272",0.0160883637144178,0.0138090510612461,0.00864777268771433,0.0199425906083033,0.00601064392811734,0.00324587532459586,0.0389235071351441,0.0203706600436935,-0.0224289272991482,-0.0175493094837592
"273",-0.0126096387278652,-0.00813448715664822,-0.00311789527239914,0.00308002919000505,-0.0102906438261211,-0.00555885636671316,-0.0155132949450089,-0.00381126965752687,-0.00279798551310539,0.0175493516543039
"274",-0.0267737316193998,-0.0500670187854794,-0.0336201815651371,-0.0538380055091345,0.00763926462169384,0.00704401338032112,-0.0316631154906964,-0.0435414723729423,-0.0159371271815292,-0.00831537447744168
"275",-0.008051893470024,0.0055215656334151,-0.0129448523459926,-0.0163761735563973,-0.00305352165609762,-0.00177668404761178,-0.019189448873313,0,0.0144844548357663,-0.00465840677163776
"276",0.00661400576446658,-0.0108826771651727,0.00573776336801601,0.0169557751738949,-0.021546541957122,-0.0112341034695836,0.0241040359187705,-0.00857177407165544,0.0101180554283773,0.0121684457745848
"277",-0.0064212474509121,-0.00353272758099421,-0.0252649012151912,-0.00188632406186073,0.0114421891722252,0.00843693240165777,-0.0310255527035753,0.00192130360746123,0.0127991321713774,0.0299014221653737
"278",0.00510991389768822,0.000911718154646524,0.0100334674308051,0.0123962256642085,0.00416215447158286,0.00223087233836239,-0.0200316208554091,0,0.00362639560439559,0.00658490632753428
"279",0.00927114815982977,0.0254022453868097,0.0149005955831762,0.0161266869160333,-0.00595164105075874,-0.00211463661948452,0.031546794441133,0.0134228940085339,-0.0218986089587516,-0.0202200517606466
"280",0.0102228058240352,0.0141137162590976,-0.00734087688391361,0.0224835215121146,-0.0105843503507229,-0.00423869837066138,0.00468076490155256,0.0085146102192073,0.00123138920337218,0.00819414455935585
"281",-0.00879947770113088,-0.00778599842136729,0.00986025982068672,-0.0128629709769462,-0.0146968990373318,-0.00548762681235082,-0.00745439279347437,-0.000938284142983692,0.00301874993249651,0.0201685945015921
"282",-0.000222043331103206,-0.00392306628506423,0.0122050357416772,0.0071343357271676,0.00767783914413678,0.00213988118937003,-0.00406842412678898,-0.00187775491620568,-0.00624230304583995,-0.00472116848927839
"283",0.00281174989695798,0.0125059915315988,0.00964661540929423,0.0130824798197509,-0.0101229042784076,-0.00719290737984513,-0.0174394485456645,0.0169331018775234,0.0272574306840732,0.0326120194826895
"284",0.00295176456185775,-0.00048654988345731,-0.0207010302620606,0.00834791206910324,0.00692722850081151,-0.000905633199416833,0.0233455420779582,-0.0129512579351064,0.0181261843606424,0.00516786232688937
"285",-0.00831370398332909,-0.00136201347290987,0.00731734818200858,-0.0140099456669825,0.0105914861331027,0.0103106520422955,-0.0226563978156941,-0.00674775112377812,0.000107271559572464,-0.00542700647917216
"286",0.00615760025028456,0.00964653537819626,0.00807102578679952,0.0134194314657685,-0.00572612107071679,-0.00280324825175249,0.0235014200835297,0.0049066603367518,0.0015013297587132,0.0137852753837973
"287",0.0126086642789431,0.0147652699882279,0.0208167857480752,0.01862334506972,-0.0102150915640399,-0.00663536466664449,0.0309277300259925,0.0140845293435012,-0.0069600707459051,0.0096317030604518
"288",0.00750061400775626,0.0194958227338011,0.01098038230012,0.0132081545501372,0.000329554876296267,0.0024902457545084,-0.000605963296015144,0.0138891589790338,0.0104593597252396,0.0213242670851113
"289",-0.00101234551709239,-0.00335833460404167,-0.00543087754719218,0.00843902086719939,0.000877936742249785,0.00237183650263706,-0.00712551960140539,0.0100455397756496,0.0114182052226892,-0.00137369983327418
"290",-0.00976670931398227,-0.00393130458355961,-0.0109203599239003,-0.0107494696568509,0.0177640861709323,0.0117172329349466,-0.0207667369199471,-0.00542502484813645,0.0127663959988014,0.0096287237141659
"291",-0.0222837780192591,-0.0247131485550178,-0.0118296197772652,-0.0397527764928246,0.0153010945047354,0.0106901587079655,-0.0174642972233614,-0.0334546569713673,0.00197939372808409,-0.0163487644500253
"292",-0.00239135762259268,0,-0.00079805824611423,0.00544369740651884,-0.00257800533374808,-0.00254170560008349,0.0053958930405329,0.00169302083010026,0.0110209814930338,0.0146813734667879
"293",-0.00382023055472591,-0.0112725307564474,-0.0231630174749682,-0.0232226880063058,-0.00971787563442272,-0.00376752172915384,-0.00805019404045382,-0.0159622122874985,-0.0211846775233376,-0.0035489822077398
"294",0.0063162689718439,0.0109138890969507,0.00572349109072445,0.0210033438310371,-0.0119699621397258,-0.00433739843600534,-0.000955159426825114,0.0160308280823311,0.0266862891363731,0.0219177486587276
"295",-0.0206979700274552,-0.011374833244097,-0.00894296760257418,-0.0342856839223376,0.00534754972563878,0.00804239701853793,-0.0458744580823079,-0.0159657780033329,-0.0124846601260268,0.00750686883795959
"296",-0.0103003538094038,-0.00887259595378231,-0.0147660370923232,-0.0138316879358137,0.00130311936317073,0.00343556377079479,0.0100169413646276,-0.0112617108925558,-0.00424874611398962,-0.0101118449885799
"297",-0.0131834453729115,-0.0102313469504068,-0.00416336097617542,-0.0175500537545958,0.0147451893725248,0.00717895914855471,-0.0161985379397347,-0.0173742609914698,-0.00228944748837334,0.0188172265118327
"298",0.0359375831858182,0.031806265514988,0.0292644355954432,0.0672569594401005,-0.00854763823200633,-0.0108565030311523,0.0710683011932141,0.0451867483106048,0.00125164281052537,0.0155672258795234
"299",-0.00935140753474173,0.00250418363338079,0,-0.0185264349540042,0.0192905756622521,0.0115287612248265,-0.0214898573963261,-0.0203008915719398,0.0106261487785426,0.0109120036113952
"300",0.00220751126084728,0.00490082020347637,0.0032494055348169,-0.00910989375559546,-0.00782405704289557,-0.00525997638028786,0.012503530305283,-0.00230252602097791,0.0137098646797265,0.00102792855388745
"301",-0.0154958900519578,-0.0253393864126886,-0.0663968792273657,-0.0354518500479746,0.0123621077658118,0.0103558723104122,-0.0163074983177226,-0.00576937859902116,0.00376248744203722,-0.00128365835410771
"302",-0.0101070265936183,-0.0171690388768914,0.0286210895299339,-0.0247063680755417,0.007684137675535,0.00501625222068292,-0.00675986764562275,-0.0348162182599996,0.00466010540634287,-0.0401027999348437
"303",0.0415432936214524,0.0303457191261616,0.0286675528931388,0.051993507098774,-0.00386530948903052,-0.00683594493682915,0.0510451047086031,0.0320642496191481,-0.0269234451330734,0.0222280619906789
"304",-0.0247697783926784,-0.0382679230349828,-0.0303275877127035,-0.0600519033094605,0.016569256805306,0.00863065584302114,-0.0109466031865481,-0.0194173655463891,-0.0358549119170984,-0.0432275970356528
"305",0.0185227310879945,0.0126927838375328,0.0185964252834616,0.0168424093909199,0.00247549157908167,0.00216560632540119,0.0417766141325915,0.00406186277260501,-0.0336414119342067,-0.0402519045767038
"306",0.0199878952862722,0.0179050834557806,0.0307055873794548,0.0383354698969915,-0.0193456879784319,-0.0176158761399283,0.0170583233002628,0.039270428680972,0.00211315750803442,0.0182596148216252
"307",0.00096505377838163,0.0177855809852951,0.0104670073118829,0.0153525524083113,0.00419804496240572,0.00352083775967915,0.00788447600366093,0.00954243526011167,0.0291898452650354,0.0100869355330777
"308",-0.01223596952926,0.00384050258767243,-0.00796820067726134,-0.00811343802672027,-0.00418049505619467,0.000767736169093647,-0.0264203077484572,-0.00378110407547416,0.0115388759342541,0.0299583839720059
"309",-0.0031531623775326,0.00124378250344637,-0.00321303627346925,-0.00483329928329834,-0.00703063135919091,-0.00131482967225749,-0.00424532191973626,0,-0.00362477600347211,0.011042175200366
"310",-0.00956461765011785,-0.00487234229195932,0.00402916849348856,-0.00179380326122958,0.0097221600871551,0.00394892107372891,-0.0153773455759098,-0.0153696568821245,-0.0169056496565979,-0.0237079151963853
"311",0.00349782995086501,0.00806374909955876,-0.00722292432046645,0.00591409148514632,0.00355859029844141,0.0017478486589444,0.00664917726495773,0.0185002196133828,-0.0159990536351454,-0.0240109860613007
"312",0.0351593878217715,0.0318065186247996,0.0291025079486005,0.0383985241808344,-0.0162751802731484,-0.00874422454105628,0.0491549981204744,0.045411653640876,-0.0392655994130915,-0.00559131338682139
"313",0.00065884433619412,0.000369075267574459,-0.00157096895453568,0.000716633334819416,0.00212987588588232,-0.00331125122886156,0.00424607545473799,-0.00271506352587858,0.0277457514650501,0.0298003766841444
"314",0.0024876495972217,0.0016609188491743,0.00472058350334259,0.0121742355850873,0.00223025221915507,0,0.0204113122911738,-0.00181456664983437,0.00168030699048871,0.0054601548488511
"315",-0.00109505221207151,0.00543389247927939,0.000783154026538169,-0.00403298502223071,0.00911598123586166,0.00764205469766299,-0.0162880640971874,0.000908984611493802,0.00928206238608942,0.00705930535222699
"316",0.000511362555996264,0.00494694799370965,0.00704225668044756,0.0132840658539539,-0.00525204581776584,-0.00659490094593818,-0.00232380193079929,0.00999054631185703,0.0101938836565099,0.0107847322711923
"317",-0.00102205363083341,-0.00911565161078509,-0.0147631125211509,-0.00546814508717575,-0.00348443716249436,0.000110473509741471,-0.0125199871965213,-0.0151078815674675,-0.0089941868815222,0.00400083423797892
"318",-0.00723613510308918,-0.00386374259821576,-0.0149841136572572,-0.0155787374285492,0.0103840720835915,0.00597460737788835,-0.0203451974248647,-0.0189914716033865,0.0214720868062444,0.0167376768781422
"319",0.00139906647275301,-0.00295541773186092,-0.00320267348738845,0.014321348574176,-0.00335541024687991,-0.00395941075573192,-0.00210658288114163,-0.00874932973793474,-0.00563445654313077,-0.0044422060963667
"320",-0.0194089203367647,-0.0163023374989669,0.00642573322021489,-0.0163073590625794,0.00673456019854846,0.00430700603466039,-0.00362002640999803,-0.0101408207576509,-0.00512143418725408,-0.00393697157603001
"321",-0.00337362378345385,0.00197738932821223,-0.00638470679764391,-0.00236877598460072,-0.0058538000737649,-0.00252948262912833,-0.00544809190654172,-0.00986545755907642,-0.00208107331606555,0.00685105097014449
"322",0.00233199538166606,0.00488694552752467,0.00722901652620522,0.0117260715031884,-0.0124065091194929,-0.00451930002736156,0.00517396177022045,0.0136046555865059,0.00603669184461975,0.0120387266780331
"323",0.0270941577570343,0.030113234305936,0.0318977856301266,0.0295786229157433,-0.00979390095118804,-0.00675511442675658,0.0431491470299168,0.0302454466802227,0.0175648366762018,0.00956836643833903
"324",0.00146119120526444,-0.0128008677391658,-0.0146828790691477,-0.00725117863229463,-0.00172074435242486,-0.00234053596667994,0.00580571179200162,-0.00422038278812442,-0.00761229787538231,-0.00461070342382686
"325",0.0104344645573708,0.0121388559075113,0.0274508255800376,0.0150956974907941,-0.000861785739724619,-0.00100611946159856,0.00101017233393041,0.00681785281051428,-0.0209593241348168,0.000514571753596815
"326",0.000505067976996454,0.00254420062722249,-0.00305326500725045,0.00507091566223616,0.00398896511624325,0.000111672239196281,-0.00994686176630122,0.00311140590769576,-0.00408301685887158,0.00128607698844219
"327",-0.00440258269704585,-0.00879093676211029,-0.0191426380429406,-0.00927299782225044,0.00343548513762104,0.000782793442157814,-0.00465929625777672,-0.00437906492617945,0.000221573407202191,0.00616493979980648
"328",-0.00159494390402637,0.00128011234584346,0.0109291190492231,0.0143842765185924,-0.00331665687796223,-0.00100566785575218,0.0115563644746097,0.00293211223155332,-0.0116317274276636,-0.00944611904816373
"329",0.004356585708015,-0.0039267186951355,-0.00772198451017303,-0.0128230846853411,-0.00848130648773704,-0.00782984927349351,0.0229937154426081,-0.00877034172319346,-0.0224164982916779,-0.0167525302708712
"330",0.00925396191280337,0.00980952519158862,0.0194551235325855,0.00735372538331847,-0.00584667281650675,-0.00135359753509123,0.00339271025707344,0.00460849515453998,0.000573217145457328,0.0183485356086419
"331",0.000215187676173567,0.000725956896574731,0.0183203271632113,-0.00191032624652776,0.00304967886565266,0.0018065472913511,0.00225388583158637,0.00642193248079814,0.00481270785422394,0.00231666710798772
"332",-0.00393893862631101,-0.00816463469936068,-0.00899518457732829,-0.0177045298650366,0.00379939547955255,0.00180261510035384,-0.0144781528939866,0.00182342760548093,-0.0214392058059254,-0.0241397522296555
"333",-0.00589635707292879,0.00301844962138209,0.0045387243295103,0.0205982040986064,0.00713942713786997,0.00315061321660015,-0.0175442508161923,0.00873477438685843,0.00978911571586338,-0.00184207728080377
"334",0.0206858716045697,0.00729540639032056,0.00903575308970539,0.0106372088748568,0.0000648413877588627,-0.000112079549007937,0.0235194611141374,0.00739690631012757,-0.0306982566486265,-0.0232005671045774
"335",0.0027633921663035,0.00153912990063376,-0.00223866480447166,0.00958044653984591,-0.0126112324447976,-0.00810074704806207,0.00170183191305728,0.0109239740530791,0.00702469358315727,0.0253710588069842
"336",-0.00480529571053645,0.000632465966605045,0.00149592719826974,-0.000735286030412841,0,0.00147448171297859,-0.00240684205698749,0.00212597260242342,0.0199810234102384,0.0207949517827233
"337",0.00866322736695735,0.00505877370284136,0.00448067257820139,0.011168249595348,-0.00720382059821123,-0.00317191064059996,0.00794865755330143,0.00212092349332527,0.00417294554907666,0.013151143431118
"338",-0.0178104379669476,-0.0171670004509912,-0.0126389235985916,-0.0297617191848609,0.00428808198816655,0.00397704139530064,-0.0294323364002594,-0.0225785526303891,-0.00935007535553778,0.00178157001672608
"339",-0.0025806103247743,0.0075902576381297,0.00451760387166833,0.0102930032753616,0.00897754489538616,0.00645085933689327,-0.000435311337323552,0.00721892932357271,0.0165462363085529,0.016260283314486
"340",-0.00186832476760823,-0.00599032647688291,-0.015741725699203,-0.0081640275609236,0.00368921630266028,0.0011243759667916,-0.00711291567968741,-0.00662975563249257,0.00206327377494908,0.015499896788278
"341",0.0112311608323281,0.0114135023851376,0.00380815349198849,0.0128573156878955,-0.00151381875893886,-0.00168432726282308,0.0213451560609883,0.0027057584908794,-0.00491878299974347,-0.0169866569386756
"342",0.000142619362755836,-0.00496527201545183,0.000758516922436892,0.00476851142217694,-0.0109354420323613,-0.00832640793510131,0.00529638367268515,-0.00845501024415551,-0.0183929076535903,0.00550965867879594
"343",0.00206399194490925,-0.00217740539100986,0.00909775205335239,0.00240609964695238,0.000438295288669677,-0.000340242937759361,0.00669202930350621,0.00598678523806306,-0.00222510835256018,-0.0161893475568939
"344",0.0125028750991436,0.0136387953676942,0.0195342197079971,0.0212723520185605,0.00908119598848445,0.00556114377569683,0.0124472529990944,0.012624301448676,0.0211267965185493,0.0113924318653231
"345",0.000912450007653387,0.0123789875322151,0.00368443206703861,0.0127329966645875,-0.00411998777152067,-0.00169308538941315,-0.00656665296049763,0.00195910124185916,0.0241379080459769,0.0145181541236565
"346",0.00273349780433518,-0.00301269783930613,-0.0014682253796966,0.000193391853545721,0.00130639278247036,0.0022611957811336,0.00759442840643776,-0.0120870138461479,0.00325478121784029,0.00148039177348736
"347",-0.00810932614033899,-0.00684319591345428,-0.00882381420275491,-0.017340530896388,0.00521937461651767,0.00304596060882423,-0.0206562417141652,-0.00791639569752955,0.0168923035786139,0.0137964968803499
"348",-0.0169144433234664,-0.00912729997061545,-0.0178039729590395,-0.0101679883212435,0.000216888085485145,-0.00236241801814607,-0.0216615749872953,-0.0126948930216672,0.0116611328567406,0.0291615105691487
"349",0.000143410287694712,0.010566024210211,0.0143504354072919,0.00291621808290232,-0.0117891529517686,-0.00653713652345711,-0.00670078317836187,0.0121232335123649,-0.0106567639262372,-0.0144037392189068
"350",-0.0134041962812451,-0.011974874380291,-0.00819050513908282,-0.0174453356779577,0.00437736669890354,0.00442471066945971,-0.00645280649455859,-0.00980020227865386,0.00274785658118737,0.00191664407877123
"351",0.00741050082655414,-0.00388913916796607,0.00300292626332488,-0.00161422063286132,-0.00675514231911656,-0.00485701351193568,0.0143176084259649,-0.00751492378172203,-0.0204976645676532,-0.0160210091301101
"352",0.00461573696355111,0.00381346745494704,-0.0112275129574287,0.0134727051604808,-0.00888621469168405,-0.00749308014212913,0.00407455880392171,0.00757182547304036,-0.00246197401004944,0.00631828367677323
"353",0.00502513729635545,-0.00597009473372501,0.0113550013825834,0.00219323937913174,-0.00719574716074267,-0.00468933095251378,0.0104350798838722,-0.00494856348014427,-0.0295041174501247,-0.0272880294777116
"354",0.00250000577591214,0.00200215008755067,0.0134730833090337,0.0034491397217804,0.00657836981697746,0.00333304275857782,-0.00401646345413575,0.00202586985260322,0.0108657378137615,0.00670297976193712
"355",-0.0103312372784649,-0.0148943041144282,0.00221567322820304,-0.0118970544050587,0.00385746366515827,0.00594213654323483,-0.0139686144593363,-0.00845537271904606,0.00583192701538926,0.0133169815653049
"356",-0.00583160042123476,-0.00295026751254479,-0.000736895308275143,-0.0180602543714575,0.0071987247876879,0.00525615453369954,0.000729704800445763,-0.0142754339255932,-0.0122783311991624,-0.023606741866913
"357",-0.00050664213463758,-0.00989345211095416,0.0117993756316535,-0.00871917640646735,-0.00890674610727671,-0.00363734149273265,0.00554621411386491,0.00921555701334786,-0.00264727219085892,-0.0149551263085738
"358",0.0199968683720066,0.0193312140269686,0.00801762356956459,0.0318167681241177,-0.0059901192616838,-0.00524763915915827,0.0251087509289627,0.00913144153086654,-0.0023081938301629,0.0379554310072467
"359",-0.0318935711916304,-0.0281265852873582,-0.0354305974891655,-0.0362303726638062,0.0129462592646479,0.00871542490239641,-0.0396429093185707,-0.0232689639961063,0.0301908743848771,0.0255972879346751
"360",0.00242100100220544,-0.00103686674217385,0.00149947264654515,-0.00255703091743131,0,-0.00716210706547749,-0.0231463215447112,-0.0138014481175283,-0.0120143726030624,0.0102211742407385
"361",-0.00497736460821097,-0.0136831399336163,-0.0217065476377354,-0.0230703521072846,-0.00650078625747308,-0.00595496742422064,0.0039238200550189,-0.0279910871925628,-0.0277303677174762,-0.00400007566573857
"362",-0.0147121775083311,-0.0154994560585876,-0.0145371121025245,-0.014963701614225,-0.00232886595963,0.00103701475371665,-0.0205954895263587,-0.00394468852001617,0.017182863219771,0.0368531702795376
"363",0.00380749102376821,-0.000874345661877496,-0.00232904526387512,0.00583171580953179,-0.0100039739198734,-0.00874619856822356,0.00614035888695152,-0.0128712928072429,-0.0163180768668609,-0.000227787839221172
"364",0.0126440902865272,0.00787889120451113,0.0101165599718052,0.0108080954858287,-0.00213358668576713,-0.00232115478033101,0.0208995086288175,0.00902690591787225,0.00268696267960178,-0.00638108513231939
"365",0.000587788544277767,0.00550056603263394,0.00924503560365464,0.00339913146498971,0.000224367096081757,0.000116687454229325,0.014345705005389,0.006958423829589,0.0137481064022347,-0.000917259715971785
"366",-0.00484463077578212,0.0012476362156506,0.006870232102411,0.00423401061545126,0.00202522244492553,0.00337321270079061,-0.0294638275962625,0.00592306152178468,0.0027582805939943,0.0101008964033154
"367",-0.00973662822078991,-0.0107362322898492,-0.0106140936308438,-0.00484892860850827,0.00842069536232604,0.00545092773367561,-0.0148755546298774,-0.0107949069039742,0.0118051461318052,0.0136363564003168
"368",0.00126594508779987,-0.00164721018015634,-0.00306496330652828,0.00155371627741197,-0.00590068168111346,-0.00576740042327317,0.0206468336573253,-0.00297625855165828,0.00158585185303406,-0.0233182687419895
"369",-0.0162313579622246,-0.0198000887288361,-0.033051837580634,-0.0326447958511973,0.00582317397987908,0.00464016402223577,-0.0247579155264256,-0.0107123795540336,0.00599410780353082,0.00688701191158803
"370",-0.000988240798294848,-0.00372095524310823,0.00715421746027078,0.00291539529866625,0.00211605611050425,-0.000461400394583422,-0.0207431121339622,-0.0207616182382869,-0.0209106358935571,0.00706784901461277
"371",-0.00197784876854634,-0.00377550485477429,-0.00789237622450323,-0.00443302921618249,0.00666599773681176,0.00531336078974132,0.000474055122355876,-0.00228624587482862,0.00436335994320181,0.000226438523680317
"372",0.00472591665324473,0.0134182353570089,0.0151877110943051,0.0200238963215336,0.000442066519066087,-0.000114998327469529,0.017652312521955,0.0177084257762081,-0.000571658847928758,-0.00384796818793998
"373",-0.0271601938061028,-0.0245603367888673,-0.0251969412208602,-0.0343104604194363,0.006729896713769,0.005630920728666,-0.0357588588332096,-0.0227224057413241,0.0364905407570473,0.0331744203459301
"374",-0.00545899761684421,0.00466271682681274,0.00565417844155558,0.00966901005454113,0.0117260086150681,0.00491330641639909,-0.00780732210606183,-0.00691275942423264,0.00949122602923258,0.00263902291314744
"375",0.00352862116863495,0.00268130985369774,0.0016066413664575,0.0075728712858012,0.000216275423075007,0.000682624967531353,-0.00327861773415461,-0.0101245600122183,-0.000765267292388017,-0.0177670229074153
"376",0.00312547275842201,-0.00874292950025712,0.00400957048697181,-0.017831006226583,-0.00236913007424389,-0.00271338506421059,0.00575669771612186,-0.010014756912224,0.0137855795670552,0.0176417854465454
"377",-0.0171366982988185,-0.015357335668614,-0.0215655204209058,-0.0285068422550631,0.00522918431561692,0.0024004735979215,-0.0207687631471161,-0.0079636975500581,0.00550392810257172,0.0190915051542797
"378",0.00103037309564069,0.00779837165568886,0.00326535179180265,-0.00285753221355767,-0.00216744135656988,0.000342217287509605,-0.0080163612298717,-0.00282077494598443,-0.0119137063843235,-0.000430672741844051
"379",-0.0102129125127394,-0.0119209909872272,0,-0.00356223885748652,0.00456247618713213,0.00467451894418414,-0.020538517789767,-0.0002172466199446,-0.00901580510570943,-0.013571687391414
"380",0.0177570173781061,0.00910147109884596,-0.00406812395270506,0.0122794598892824,0.00648718925110692,0.00249699759628386,0.0723616036747416,-0.00217642184936562,-0.00405570522671139,-0.0362524577358925
"381",-0.0192548939324572,-0.00985841907785334,-0.0163400688547592,-0.0201917990952445,0.00440394052384119,0.00475399320032399,-0.07356963870567,-0.00719771392295954,0.00704379257050647,-0.000679765429519197
"382",0.00408694155240208,0.00646121536363364,0.00913612776745265,0.0181009129705274,-0.000107367202276887,0.000338498289032652,0.0181663330653778,0.00395456803721594,0.0221857814207651,0.0272107961405996
"383",-0.0116523372741529,-0.0181014693275593,-0.0131687109344015,-0.00669624794779611,-0.0142259832414862,-0.00934835704377379,0.000339831593961559,-0.0205692975039501,0.0174276169937733,0.0139072576091852
"384",-0.0090434283978641,-0.00321542593869406,0.00667222000372059,-0.0012396896267165,0.00878959424145687,0.00534350321173482,-0.0348223051038647,-0.00379771828928366,0.00788146246820243,0.000435523166912199
"385",-0.0140976291743878,-0.0148387082721269,-0.0165698420931774,-0.0166798209970431,-0.000323236190593823,0.00361806671899312,-0.00950388107791444,-0.0222020872242593,0.00271081210673296,-0.0317736170793276
"386",0.0245477872725828,0.0128792369208048,0.0252734658336937,0.028875990562206,-0.0180758195052192,-0.00912654168660398,0.0701849078878423,0.0155958033286954,-0.0179889366328155,-0.015284340931413
"387",0.0100029494938407,0.0223062152833959,-0.00493012718655683,0.00467730756450924,-0.00515072959657781,-0.00477573938168707,0.0161046345704441,0.021906593246759,-0.00232953192864194,-0.0235107378302527
"388",0.00623067121954768,0.00980263063852416,-0.00412879067245309,-0.00862447775960651,-0.00374483262948266,-0.00342785680208391,0.000327070205614399,0.00773467129290895,-0.000530704727969455,-0.0170640232062798
"389",0.000555265089721368,0.00584585172897589,0,0.0123954266068698,0.00386977141297784,0.00229321401638072,0.00294015991922847,0.0164470297507491,0.0100881917826949,0.0121285500252375
"390",0.0113448771856073,-0.000104032210217819,0.013267459255667,0.000608010072664422,-0.00495581478061746,-0.00343108479443666,0.0317590875911817,0.00539379651034722,-0.0216569063817208,-0.0218516034181685
"391",0.00541239230419532,0.00352893647607755,0.00654636549939802,0.00144407686223769,-0.00199266027200573,-0.00160758532293603,0.0213098773972331,0.0313306908640267,-0.0267569100957857,-0.0225799169704837
"392",-0.0207536890585488,-0.0212016744894962,-0.000813031652907581,-0.0369584911084186,0.00975903589449545,0.00862301067035909,-0.0615145624632232,-0.00728271180086204,0.00839132162967871,0.000737439518115224
"393",-0.000239082649505118,0.00612833729991769,-0.0113914361617979,0.00685556738653337,-0.00999405394295594,-0.00581380419161526,0.0151515634700914,-0.0253612858592421,0.00394174961257554,-0.0125246920014604
"394",-0.0146638899977006,-0.0149128282375967,-0.0115227950903365,-0.0169050685350693,0.0100949433513606,0.00573308787685378,-0.0212526464263304,-0.0109678782721471,0.000436263487048283,0.00497402307860817
"395",0.0213525589425771,0.0110874892033701,0.00582884639947867,0.0554093889836158,-0.00406313378914891,-0.00285020347145815,0.0500583703878972,0.00217452948492869,-0.0124278530765991,-0.0113834159100783
"396",0.0178176080603243,0.00991134202375621,0.00910562598235742,-0.0104094701863132,0.000992430824902524,0.00194396665113428,-0.00489359182435345,0.0197439537019786,-0.0118114477011346,0.0197747231077408
"397",-0.0132263044341787,-0.0110669628345497,-0.0155863847070056,-0.0224103155585547,0.00991492183246812,0.00798691539106011,-0.0117386787247815,-0.00531931965053034,0.00625564140713708,-0.00834558517007378
"398",-0.00528281072684766,-0.013091238983021,-0.0141665766963927,-0.00678376046675078,0.00221171250181373,0.000499198946139146,0.00240778790115281,-0.0034221626674299,-0.00566165617980341,-0.0111386394825681
"399",-0.00927397293500165,-0.00363737086224336,-0.0253592271586777,-0.0306166557357118,-0.00229395355297723,-0.000681037598829093,-0.0140912721690194,-0.0223228465330827,-0.0159651780730155,-0.0330412197272842
"400",0.0269622667555269,0.0300623911798867,0.0225498955672205,0.0128764643056065,-0.00744545473037894,-0.00511197850344747,0.0427156780025122,0.0208565725678271,-0.0233718745560686,-0.00698947251736459
"401",0.00444035782124708,0.00145922019301037,-0.00593722783683248,0.019909105669907,-0.00408227011098494,0.000342157095583051,-0.0046728586410032,0.00559124024448865,0.00650554120572644,-0.0106882484373897
"402",-0.0148918122491363,-0.0185263148524168,-0.0221842992481058,-0.0343371034935692,0.0162836075404598,0.00936069364257097,-0.0242568840360757,-0.024807436540324,-0.00634814180918908,0.00553359520466379
"403",0.0185813757699709,0.000424413835264259,0.0148340046112698,0.00243565677023416,0.00272409970330245,-0.000452422573219757,0.0323977213618298,0.00197367000077353,-0.0192821010236776,-0.0280398631922217
"404",0.0103582019033113,-0.00190784419451351,0.00601878141993506,-0.0104472810479204,-0.00956476624979163,-0.00486553247093868,0.0245456260195087,0.00656592726293126,-0.0390856686012081,-0.00107836893611957
"405",-0.0104047274027457,-0.00488557886218177,-0.00683767787493084,-0.00834759934866391,0.00932840590874817,0.00693576771036919,-0.0221378278005669,-0.00478363728496045,-0.00751879727050897,-0.00863694178083629
"406",-0.00603032559218808,-0.0175027824351039,-0.0172114575644197,-0.000247602862745722,-0.00347924356568285,-0.00214516221419636,-0.0161266652393151,-0.0190076739534224,0.0129160586034298,0.0334875668411299
"407",0.00754438281673431,-0.00695175527801906,-0.00612948555996273,0.0131250378865178,0.00643720103016787,0.00305581389444076,0.016548783784762,-0.0144768315541705,-0.0270966166526879,-0.00869334665424149
"408",0.00486320012741737,-0.00700066669352362,-0.00704876746058025,-0.0156437982757692,0.00867340032354869,0.00372310562816747,-0.00155058962401089,-0.00339020285381186,-0.0216761316112446,-0.0135530788405448
"409",-0.0136740690578961,-0.00638938226601327,0.00887345331524769,-0.0168857787720098,0.00397653863615011,0.00247226884589358,-0.0209626359133895,-0.0068027449089586,0.0150715708516644,0.00565732592459312
"410",-0.0109046145090913,-0.0121949587640928,-0.0158312478138131,-0.00833590629245962,-0.00385416069721634,-0.00145790323890693,-0.0206187835656048,-0.0228309300775357,0.0206852403292421,0.0155371930081818
"411",0.00464630258543197,0.00224490547322698,0.010723902753645,0.0254714332614916,0.00279467698042857,0.00291940065353291,0.00242931165175242,0.016355034505432,-0.00460029839612097,0.00791332262534139
"412",0.00172437858738195,0.00515096446918339,0.00618888754352098,-0.00149003563515548,-0.00182212297054396,-0.0021264685954494,-0.0137316265725805,-0.0114943220406781,0.0279790788903094,0.0429208050077479
"413",0.0144756676741828,0.00713019897673517,-0.00702966029167174,-0.00074672994406666,-0.000644244946379047,-0.00291732652079113,0.0229317862840279,0.00907021593364354,-0.0148238269201523,-0.0338770128588113
"414",-0.0202855646221695,-0.016371873923633,-0.00884938912388411,-0.0206621075101745,0.00999180153880341,0.0066385650066636,-0.0220979534492141,0.00230478698580061,-0.00185004928835575,-0.00571443886543999
"415",0.00291308420444647,0.00382387204602463,0.00535692202382987,0.00177973885539418,0.000850853208089974,0.000335705926067575,0.00769630166842261,-0.0043690429203106,0.00370694427282814,0.000522586882356402
"416",0.00973399699532473,0.0109791295106587,0.00444065309947428,0.0213139927026871,0.00170036485103209,0.00145289831660422,0.00893753343029347,0.00808308739197283,0.00160036926257412,0.00939941240979691
"417",0.0121276308168037,0.0141845439877004,0.0079571525073765,0.00695658502181407,0.000105782307984637,-0.00145079046557905,0.0331773659485071,0.0119128681418854,0.0100786503186008,-0.0196584834087645
"418",-0.0107534031544112,-0.00611898968346025,0.000877324077001695,-0.0118431951460081,-0.00445508194181687,-0.00122939918409826,-0.0112240076940676,0.00271665735732185,-0.00571916524701888,-0.00369406808285622
"419",-0.00621192650062152,-0.0127529203571466,-0.0131462464845543,-0.0302120728212184,0.00930392423206694,0.00544423363304958,0.0122971971154322,-0.0054184666923428,-0.0307184191741331,-0.0259532462648115
"420",-0.000859086133995213,-0.00467697943394185,0.00444065309947428,-0.0164777676458648,0.00423939141187701,0.00245640848100748,0.0137049329474175,-0.00726426690777138,-0.00391411630987804,-0.00570970809837212
"421",-0.0301063228249987,-0.0449765390571768,-0.031830468761617,-0.0460733661184207,0.00801951824575919,0.00501122648440955,-0.0311871724281207,-0.0420764719756538,-0.00633793898260793,-0.0142191914588167
"422",0.00314426237804932,-0.00562320196070454,0,0.0142699915289932,-0.000524442836401184,-0.00221559428934992,0.00634302807327791,0.00501258281870154,0.00752652133596787,-0.00998620532375682
"423",0.020655680691289,0.0172008771741994,0.0246577594428641,0.0124460117889942,0.00419021049638912,0.000110605937233776,0.0431770592124003,0.0261287020835204,-0.00151939725806294,-0.00224151519185878
"424",-0.0296870856994478,-0.0277971033402328,-0.0276293905549236,-0.056119898025603,0.00990814841019638,0.00455298961216477,-0.0438067460694841,-0.0199074117666342,-0.0300532966008965,-0.0365066424621719
"425",0.00405765407844982,0.00428871248294138,0.0128324446561443,0.0161382924211084,-0.00619598768696294,-0.00254308511241186,0.00537087651286905,0.0243264574509607,-0.0296770435266582,0.00145725716199618
"426",0.014468133394469,0.00142334361628205,-0.00542974949048536,-0.014767321253086,-0.000520174353783598,-0.00177285502768076,0.0114708699775952,-0.00806978307659911,-0.0153597276292141,-0.00844003600158705
"427",0.00462114395182267,0.0234544059271871,0.00636941891916298,0.0333708636673198,-0.0128919923963501,-0.00499564997812285,0.0105639702084996,0.0167361932402896,0.0337985896606847,0.00675078805886775
"428",-0.0475850529336085,-0.0467593354223661,-0.028028898843431,-0.0785440887403678,0.0324408349204721,0.0191917000490742,-0.0614908289731306,-0.0477823497888562,0.026604830181145,-0.0393584528508193
"429",0.0167374580722355,-0.0118991489022418,-0.00930256531601337,0.00861295377684623,-0.000204342020202808,-0.0028457514324115,0.0307943062381089,-0.0177670625292086,-0.00992775941020507,-0.020333922337049
"430",-0.0449631340170598,-0.045956821531111,-0.0356806867531775,-0.0709656663581808,0.00500027104659573,0.00900235036394115,-0.0465598970389414,-0.0381322933197102,0.11290529869898,0.0300495994542949
"431",0.0296715227281901,0.0569291114278545,0.044790691650513,0.0843105905407147,-0.0146204203859125,-0.0117521777720602,0.0845004182413953,0.020076247261424,-0.0311256263880836,0.0018046140202741
"432",0.0397139456533044,0.0714108626885557,0.0540540495153572,0.124525141411412,-0.0317368580044692,-0.0178372096392191,0.0327336483931435,0.0652989844072287,0.0384057957099349,0.0330228692629901
"433",-0.0226394744464377,-0.02047301328105,-0.0344826139508997,-0.0652458467083256,-0.000105608296371962,-0.00212933853845132,-0.0880951386994837,-0.0179793836952259,0.0372179214741364,0.0345829335306627
"434",-0.0227518798907062,-0.0234552950217517,-0.00915796510052336,-0.0311455414726306,-0.00383211337374612,0,0.0063640050325191,-0.0158998814764973,-0.00964341780668332,-0.00983125370641769
"435",0.00320581073466175,-0.00190264994680089,0.0138634271540574,0.0114812158670423,0.00438108940303583,0.0025835119674118,-0.00739028894017635,-0.00612003643640513,-0.0182291779891304,-0.00822696864585204
"436",0.0156394454073692,0.0243029610423737,0.0173200828746365,0.051361710393625,-0.00202191846885891,-0.00302642479536919,0.0185311653390003,0.0187189280874203,-0.00299852384959665,0.0174484640515546
"437",0.000496608543807175,-0.00930442167165191,-0.00537652638102559,-0.0340080471130192,0.00724849507256309,-0.000673455086094621,0.0207925776335842,0.00580278741375828,0.00219782540883151,-0.0118076703580804
"438",-0.0783618224020873,-0.103545580552664,-0.0774774041102719,-0.116792218785436,0.029100437360839,0.0139463479056081,-0.0598349294205924,-0.0973557861729982,0.0338181098086114,-0.0620198269049511
"439",0.0413899883106008,0.0440025160970077,0.0410156415542433,0.0809867363154271,-0.0243699984445532,-0.0132002378979045,0.0485783586324779,0.0162451331775211,-0.0502400357262476,0.0279040396033075
"440",0.000603506902418172,-0.00125489258822475,-0.0121953064462307,0.011999126103444,0.0125804297298446,0.00704951037214019,-0.01533464445627,0.00943394339526638,0.0105795345009991,-0.0233106248146986
"441",-0.0362741310484452,-0.0419492621312614,-0.0427348635694603,-0.0876230412326523,0.0080392430364693,0.00560094178108939,-0.0662296572099632,-0.0501039442464298,-0.0423403391608662,-0.0552870733393158
"442",-0.0135001831017242,0.00209777872987749,-0.0198413087382803,-0.0263073843568067,0.00880372802830776,0.00378716130252799,-0.0533707113227451,-0.0213173616136897,0.00315794963784888,-0.023345023034933
"443",-0.0509337511473518,-0.0580848254138944,-0.0323886010824155,-0.0751952906139518,0.0181724926749822,0.00809961518085545,-0.0183605825642333,-0.0823793950792684,0.0204625630445605,-0.0425672076916122
"444",-0.044785757007434,-0.0500000664301598,-0.036610776729827,-0.0777897827809801,-0.00302525051080271,-0.000770303335253519,-0.0844509329595455,-0.00182558530757593,0.0354769581807897,0.0123118879564208
"445",-0.0251927597930937,-0.0102340295612176,-0.0369163518871155,0,-0.0143619316698953,-0.0127777980928813,-0.0167153224577167,-0.0423782018800829,0.0246361988530834,0.014527083835969
"446",-0.0698387243329397,-0.0747412056207259,-0.0462234727307558,-0.0736638589607006,-0.00841533651539106,-0.0100432205854216,-0.071563087075935,-0.0799108206213267,0.00536797149111989,-0.0466200320130208
"447",-0.0242560663222771,-0.0249042994859816,-0.0437350761719814,0.0115369272216319,-0.00703602253460522,-0.0117221607954376,0.0795657164041759,-0.0311420042491198,-0.074304792562741,-0.0443590389076348
"448",0.145197740708131,0.137524656236034,0.158219997006472,0.227698445648615,-0.0128197815244123,-0.0068427865690569,0.0747488891864938,0.10714274079544,-0.0147801368086982,0.0555555194676047
"449",-0.0148002152361718,-0.0184228360656959,-0.00533610937857576,-0.04976776000617,-0.00643989050073412,-0.00470789581773434,-0.0648742517252026,0.0438712978247984,0.00256127582781485,-0.0183518618979334
"450",-0.0984476316246472,-0.105571671603791,-0.104077325824267,-0.161661996368433,0.00956327774355081,0.00819154695801338,-0.141666865547044,-0.0908530182383238,0.0135036622933209,-0.0455026021484503
"451",0.0416571578762153,0.0498359307126894,0.0610777784091849,0.0491463003845827,-0.00515797901341142,0.000229640606186798,0.0628644157843998,0.0472466334707715,-0.0482534761314001,-0.0188469788539656
"452",-0.00597191088290949,-0.0162398209509261,-0.0135440042860739,-0.0313616605974704,-0.00687671031564752,0.00629255115264571,-0.0102766263022904,-0.0327814998882823,-0.0262328411371821,0.0112994087772322
"453",0.0600796186373747,0.0520634726687559,0.0789475275682674,0.0700818275274318,0.00799021861925375,0.00102330629204883,0.00946015358184771,0.0620804816764222,0.0167076935203692,0.0201117479402557
"454",-0.0298553081930782,-0.0585395313191984,-0.0360551962160827,-0.0796631243989907,0.00528412762720243,0.0105631926281442,-0.0345142305126829,-0.0423379036707764,-0.0314649808917197,-0.0357795082209367
"455",-0.0544544043277595,-0.0762821322098519,-0.0605061147916494,-0.105284992279647,0.0202904169477158,0.00764337054877773,-0.0733901208563129,-0.0514682512166612,-0.0568196771908416,-0.0473305935845669
"456",0.0115841783422352,0.0183900955359495,0.0339579502725404,0.0279071627819261,0.00741907053811408,0.00133798296734344,-0.0155853317146696,-0.0285216673763252,-0.0147817182370898,0.00397460927152582
"457",-0.0507144694542776,-0.0494037030429747,-0.0600226146588918,-0.103167699046605,-0.0106376710448732,-0.00423253326698969,-0.0641057244124386,-0.0748297170577805,0.022080636317604,-0.0399841171555951
"458",-0.0355009651348255,-0.0580644979122779,-0.0602411090229161,-0.0262359274257586,0.000723673204495512,-0.000559311287050668,-0.0521350538779515,-0.017027996708558,-0.000415441080396484,-0.00742275787031688
"459",0.116855471311958,0.129756407405619,0.12179501469768,0.209326374468313,-0.0145661908229018,-0.00805915290467119,0.163253182144635,0.0362205735460992,0.0223053615960098,0.0274200670797233
"460",-0.00725271549552642,0.0148197449463972,-0.0228572534722251,-0.0317052614484162,-0.00503114016540518,0.00146640935882969,-0.0397386891146865,0.0136776423621587,0.00284590048995925,0.059037684233568
"461",0.0345941039693194,0.0288751588378855,0.0538011128977984,0.134956226106578,-0.00906165609680964,-0.00766110052027713,0.0484548269650786,0.0468515451841667,-0.017432445945946,-0.0412371829495353
"462",0.00550350542809408,0.0125803927063963,-0.00110991013524375,-0.00857742969687492,-0.0129717553705626,-0.0020442670280556,0.0629526469872164,0.0204080925337844,-0.0188420164879936,0.0111509323669647
"463",0.0028915934646907,-0.00382289084457454,0.00666662684671815,-0.00904420231376379,0.00270338711691709,0.00159840793000376,-0.0364277047636143,0.0245615343736463,-0.00336414372661309,-0.0110279603272104
"464",0.0339821481535669,0.0697155567244283,0.0551877856336327,0.0912697328553296,0.0187686299540744,0.0119714229517294,0.0556098560339779,0.0352741715220719,0.0616034475837819,0.0454003257497158
"465",-0.0420274993404275,-0.0594918678766143,-0.0209206682314618,-0.12727269115983,0.0118575247745756,0.00529535511538359,-0.0965803155190601,-0.0370490679093639,-0.0355060929184117,-0.0259048539988933
"466",-0.0554113067673299,-0.0632549829067478,-0.0865383196228724,-0.0504167558267562,-0.00721938268540423,-0.00302650654899261,-0.0452688146275562,-0.0398495457345551,-0.00796706011124759,-0.0438013163797875
"467",0.0330177451636124,0.0563285900453008,0.0584796812905737,0.0811759562980416,-0.00653446027009341,-0.00359710817738434,0.0592021179806264,0.0296964933025841,0.00387702847027116,0.00122699958366002
"468",-0.0131042525475108,-0.0215225576736183,0.00883963570798674,0.00933438012124377,0.0048795111188249,0.00101555596279446,-0.0857360737628258,-0.0535096962064453,0.0148965793103448,0.00653592119552315
"469",-0.0308759346219815,-0.0252792140786825,-0.0416209199757402,-0.062323983893002,0.00295604005116479,0.00371907856173137,-0.0127251835296606,-0.032672537045115,-0.0207936797827213,-0.0190745666179768
"470",-0.0440011701248243,-0.0565846788451937,-0.0274286767090256,-0.0741851130280218,0.00642181871995118,0.00617626018073403,-0.0736898414709209,-0.0288424985236464,-0.0284525040200208,-0.0293754072624588
"471",0.062339512076196,0.0828275129396723,0.0681551806375833,0.138489720477353,-0.0239525540882518,-0.00725445096683863,0.110708085292271,0.0441579256230675,0.0307143142857143,0.0187553871036426
"472",-0.0499067987144763,-0.0524233593732462,-0.0539051978339044,-0.0960128352126198,0.0198246966408915,0.0098918942156323,-0.0985839050653171,-0.0550149001300444,0.0159390293571995,-0.00627609242624128
"473",-0.0132757924835234,-0.0327068421421542,-0.00232582275416837,-0.0166515374284436,0.00441321883027612,0.00423015778316826,-0.00785495431997674,-0.021386170030963,-0.0088676804010499,-0.0227369028419511
"474",0.0188368349593959,0.0143883829064757,0,-0.0146453125163503,0.012867757937171,0.00775920959401577,-0.0401949375588376,-0.0129503731629449,-0.00192704743490579,-0.0150796573222827
"475",-0.0640789845033101,-0.0606381305984661,-0.0641026345555075,-0.0863913876468111,0.0256149810331636,0.0107787950316738,-0.120558514761952,-0.0873306021825038,-0.00344780020830782,-0.0113736460813515
"476",-0.0742332061131772,-0.0683277717170022,-0.0286425613635201,-0.0716825430733999,0.0516613557736054,0.0201301840622463,-0.0873017501618832,-0.0336927773725539,0.016468239234203,-0.050884855047417
"477",0.0539427766187364,0.0571312878026542,0.06153835906308,0.144030280645251,-0.0144595861402277,-0.0091733341873258,0.0826087906899478,0.0418409190886899,0.0735194175705685,0.0172494312916369
"478",0.0692910456326812,0.0770407414171292,0.0471015499385763,0.0607947693653297,-0.0156431334974173,-0.00936599135575567,0.144578491181861,0.0441768282603312,0.0261256316074987,0.0687441540990277
"479",0.00740933315038594,0.0202850789638482,-0.00461374391067959,-0.0189530970977361,0.0294141036869937,0.0171694225716563,0.0271133039566225,0.0209402204402886,-0.000494388802650403,-0.0334477063449429
"480",0.0386408023005822,0.0177885206549762,0.0185401688462636,0.076357410575459,0.00134301523049363,0.00609134334615047,0.0456520118736892,0.0397657288981035,-0.00605918117747561,0.0319432230558587
"481",0.0125882962396675,0.00342697951998283,-0.014789517391351,-0.0192310928479835,0.0123532089807168,0.00201714785974172,-0.00861276931710253,0.036231502831606,-0.000870850990452365,-0.0434221329352545
"482",-0.0885779266399073,-0.0877732754852889,-0.0577368645551929,-0.0962960888415745,0.0382946008097482,0.013535172436173,-0.2061117855679,-0.0784768344829457,-0.0580251041719612,-0.0310112387636797
"483",0.0384846766265761,0.0490450752943785,0.0502449395488471,0.0631625326994416,0.00383997421060922,0.00524597312738373,0.137736154270732,0.0408936074165973,0.017184335302463,0.000463807880641598
"484",0.0240419533036609,0.00749466893474793,0.00933502179619028,0.00816359120127208,0.00282217834554599,0.00156495896676501,0.045439578496933,-0.00648046913376021,-0.0100064591295564,-0.0115902577741106
"485",-0.0231334294783792,-0.0262129126797351,-0.0393061479411184,-0.0427352556716691,0.0197034978831407,0.00625241487665162,-0.0164974983807036,-0.0342437944766737,-0.00892622735626158,-0.052532722436711
"486",0.0308322068738727,0.01527811808072,0.0156436399985977,0.0592107949307461,-0.0162060251451537,-0.0105621559890778,0.0964515237714711,0.00253270948208995,-0.0129801721854305,-0.0247524516760373
"487",0.0349139392048536,0.0458618179222869,0.0450238653208814,0.0638860778518957,-0.00217260036490186,-0.003768017860872,0.0941448229702742,0.0484208968588495,0.0225442843214285,0.0461928228227908
"488",-0.0164834271824134,-0.00548143325269823,-0.00680274726266294,-0.0137613988815016,0.0197749512709411,0.00850967472386954,-0.0717928047743559,-0.000803086867952274,0.00170610242937408,-0.0218341123036047
"489",0.00681558624070777,0.0285910737315715,0.0216891303500444,0.0596194254945301,-0.00240115826406462,-0.000936850664771671,0.0663381811397488,0.0478297057136525,0.0448054226436416,0.0302580101527612
"490",-0.0240814671388502,-0.000669787504884778,-0.00335175138975974,-0.0255384687907962,0.00196132903276358,0.00604659821329578,-0.144254328055658,-0.00460291149986691,0.0112852915360502,0.0317765472120874
"491",0.0119397295004107,0.00502670244152359,0.0224214017681394,0.0139231260509343,0,0.00279872081548294,0.0946031816097859,0.00346845207897672,0.00198383132092173,0.0219319417556862
"492",-0.0139341433519257,-0.00200079329995517,-0.00548228679836626,-0.0133282865355361,0.0113913833631323,0.00216950974775232,-0.0284223876550673,0.0145924239753177,0.0221507244685244,-0.0282931297013179
"493",0.0470658289192607,0.0648182050198605,0.0507168280111758,0.0798200227428358,0.024724112615393,0.0158818188434726,0.121791230315622,0.0264953610060139,0.0225181724580672,0.0143198584309669
"494",-0.00968671596328485,-0.00972714357631699,-0.00209879093809884,-0.0174373372552186,0.0271345497386981,0.00680129185418821,0.0252791075722243,-0.0092183501845976,0.0114847384736532,-0.0136472101417828
"495",-0.0186833434827568,-0.0323192488455438,-0.0347003424541275,-0.0219907620676691,0.0209824590146159,0.00675504662555837,-0.0788995013857503,0.00446607679221733,-0.0182605290881425,-0.015267213431192
"496",-0.00430198459125108,-0.0216109358116564,-0.00435713048409592,0.00355023608360927,0.00106501016213323,-0.00330452250196855,0.0495914255007119,-0.00156787454575813,-0.0147848569887377,-0.00678285373721177
"497",-0.0128128302991199,-0.000576073234180963,-0.00218850979457197,-0.0373427066872677,-0.00768904146402094,-0.00261299288995942,-0.020939606345632,-0.0332707994133965,0.0100448024946678,-0.0282925977976181
"498",-0.0103377155993962,-0.00576480657565559,-0.0171363077248726,-0.0082815737137395,-0.00131872143971112,-0.000503874275916139,-0.00759252804603916,0.0228151513339083,-0.0099449078593925,0.00401600906206068
"499",0.00580312169796326,0.0133013559389972,0.0123734019132649,0.00709816834233767,-0.00214575055145949,-0.00100735642718308,0.00765061555924218,-0.00189058830614441,0.0100448024946678,-0.0154999422095188
"500",0.0057697551378364,0.00807837550437251,0.0188889768460672,-0.00331662487821793,0.00330857246586036,0.00534703547030269,0.0132175279106479,-0.00378777883106629,0.0256410139664631,0.0157439728792961
"501",-0.00286809861888027,0.000333731522892844,0.00763355580142022,-0.00166403916327851,-0.0011995110263574,0.00220600430128637,-0.056342164449801,0.0112015864692563,0.00876168244770281,0.0110000038080995
"502",0.0237022013722448,0.028371116031616,0.0281384433655503,0.0266664474590708,0.00952422696690181,0.00140721606045502,0.0452939518012083,0.0113038105630268,-0.00521130295799199,0.00593463684071205
"503",0.0142748081192003,0.0107108726298064,0.00842108101380035,0.0133929667593877,-0.0209191736766087,-0.0110404558681261,0.0475522128583235,0.00894186018229726,0.00721763661891428,0.0417896661742048
"504",0.0301415817166073,0.0105970979289924,0.00521930962369654,0.0476571585314918,-0.0251363207855503,-0.0143108975506198,-0.0273971537016581,0.0347121918797981,-0.00335175693545164,0.0349221404623925
"505",-0.00118355629583111,-0.00953269834100368,-0.0249221681943944,0.0129968861791459,-0.025783707060185,-0.00174999832375644,-0.0196081776772674,-0.0071381161873052,-0.0202945603515751,0.0104879131647666
"506",0.00667757498619515,0.0121912254820056,-0.00958510050571726,0.0226417027888552,-0.0100574104947569,-0.00061909617836764,0.0495778654725381,0.0273187136638842,0.00769405749192509,0.0261732517063458
"507",-0.0299558978752289,-0.0117276266568577,-0.00967696705501819,-0.057564631112096,0.0039206855062428,0.000206617446420365,-0.0338168527878818,-0.012946175745239,-0.0279572076103797,-0.0510114152463199
"508",0.00408083282072957,0.0128290300718974,0.0141151304244,-0.00430705309002799,-0.000798911606802788,0.00268298372677855,-0.00444424720384706,0,0.0206646404833837,0.0037070854943253
"509",-0.0214193927555595,-0.0345159147313906,-0.0171308039913455,-0.0216278783731019,0.0015107209566223,0.00463083071816972,-0.0460381080006529,-0.0212691420938745,-0.00639357099684534,-0.0115419980752803
"510",-0.0240208448494063,-0.0272216311773992,-0.0119824577068351,-0.0422027997553172,0.0103786483469352,0.00624872969068746,-0.0582035737645157,-0.0315100623423267,-0.0376548626705163,-0.0453058901349086
"511",0.00184070872467035,-0.0188806430727988,-0.0187429987589545,0.00293757440194975,0.00105369962469881,0.000712882544757321,0.0301237046210372,-0.0373972379219601,0.00148582215240656,0.0166340748254159
"512",-0.0314546895141599,-0.0474229712737344,-0.029213626711862,-0.0485353209136814,0.0164880599697861,0.00559511786288436,-0.0518539595104438,-0.0470086165090017,-0.0134767067313318,-0.0139557828393829
"513",0.000355626609123139,0.00649363763934363,0.0127314981993796,0.0114333867319569,0.00164001257891622,-0.000809925717414006,0.0289347253640648,0.00163030224116567,0.00751971415566222,-0.000976072559683128
"514",0.00781965666677675,0.0014336596681257,0.00685738693227522,0.0108694847090567,-0.015420013595718,-0.00921312711861022,0.0367737033851432,0.00488422198528116,0.0288593112185509,0.00439661793669699
"515",-0.0527860936317063,-0.0776664697728162,-0.0431330212158881,-0.0744086215690403,-0.000174688294181213,-0.0015320901010023,-0.108196248853586,-0.081004503163104,0.0218836660849193,-0.0311282811770387
"516",0.0431924642621846,0.0364762755370478,0.0438911438324963,0.0543684427607871,-0.0315891399760623,-0.00890448761967477,0.0995986189815377,0.0599380545581201,-0.00437760308959789,0.00401600906206068
"517",-0.0154671430371517,-0.024335008932774,-0.0250002284631201,-0.033054727333845,-0.0192466972993066,-0.00660911325139546,-0.0507600200424264,0.011226976826499,0.00510992263553356,-0.0129999764309525
"518",0.00435055113258231,-0.00652335388624437,-0.00233085376371234,0.0127620600759768,-0.00783042738723283,0.000208099472754242,0.0317003305504215,-0.0143913940838877,0.0467013112626791,0.0466058108368732
"519",0.0068581107043848,0.026651245473311,-0.00116821925861665,0.0117014676118894,-0.00872939124370931,-0.00249414125868552,-0.00838011212373513,0.0070923895524273,0.004744131986266,0.00193618162824372
"520",0.0101580182129184,0.0161772767708959,0.0315787761217261,0.0177937071367347,0.023513152234268,0.00656358008397828,0.0181536679308798,0.00289915942634367,-0.0064080946512004,-0.0270532163348416
"521",0.0338337437473089,0.0373935852287932,0.0181406155281416,0.0506994194776456,-0.0249859649007327,-0.00641701876867273,0.079618689301306,0.0177614811730722,-0.0108621750688677,0.0238332003545942
"522",-0.032497588132304,-0.0456815776461882,-0.0378619893120893,-0.0507488176234754,-0.0229985872477937,-0.0130228888990417,-0.0783031342994708,-0.0300326872594531,0.0237932057605399,-0.0121241352363949
"523",-0.0203431240252913,-0.00710567735173007,-0.0243055247930273,-0.0074498191118928,-0.00317051442263827,-0.000421918720398429,-0.0318191971026548,-0.0121334603478929,0.020223441340782,-0.00589103658931234
"524",-0.00301827207401306,-0.0128057682545287,0,-0.0101546429267457,0.0186056537815473,0.00811210457750433,0.00638118766080553,-0.00465939781653313,-0.0270507288807519,-0.0192592500730235
"525",0.0140469366979814,0.0335750123350051,0.0189800381224619,0.0298842576891964,-0.0238168926180726,-0.00861338812991019,-0.00380467024505993,0.0144684009338878,-0.00416473454141086,-0.0115811681446749
"526",-0.00489627817972982,-0.00996687366650839,0.00931307979201668,0.00736259793953797,-0.00349902403975277,-0.00508623112891926,-0.0235518623661718,-0.0151006411599683,0.00802530792330391,0.00560380148302553
"527",0.0148807958107318,0.0193885996573422,-0.00346036464184596,0.0210660074660363,0.000877911960352806,0.00234288888922363,-0.0153191229090188,0.000425762620492431,0.0105405135680645,0.0222897741548633
"528",0.028497381036555,0.0263350578528203,0.00578704777000749,0.0501052328453058,-0.00311845990165538,-0.00605609680923858,0.0685201760424734,0.0400169792935521,-0.00588112497066828,0.00743300010297254
"529",0.00137924641596343,0.00819669777487153,-0.0184119263258345,-0.00521241543404549,0.00322549892061286,-0.00203115922200137,0.0136308877698055,0.0122801875268115,-0.0141756452361044,-0.00541064938474589
"530",-0.0458091600615479,-0.0516085325172126,-0.0351699818089071,-0.0604593446435894,0.021730954530317,0.0133888227909869,-0.0858802426703438,-0.0477154022562688,0.0213994451992754,-0.0128586343260043
"531",0.0058956313698888,0.00782718261760618,0.00486042803947395,0.030029651126112,0.0129710318226974,0.00771572919398777,0.0254096126332239,0.00127380455044301,0.0230573331455197,-0.00601204533501087
"532",0.000717684682128628,-0.00517763000793647,-0.00120936469438793,-0.00624695519560892,-0.00941503327669069,-0.000314248830991071,-0.0146722905465662,-0.00296871617571792,0.00953512829629299,0.00151228372584122
"533",-0.0107577289509744,-0.0115239713187402,-0.0266344163556357,0.00502899046873662,-0.0266134707573712,-0.00786883582710152,-0.0598943124015048,-0.0110589210894402,-0.00665444899977352,-0.018117878429032
"534",-0.0427744695912257,-0.0590450852134708,-0.0335823219179268,-0.0638032380987205,0.0311488387694097,0.0168147811202004,-0.0630060273863847,-0.0692473067107666,0.03133434798484,-0.0558688131967552
"535",-0.00239833789862898,-0.0043962328474294,0.0077222844901228,-0.00712673854055212,-0.0085224870138757,-0.00728003554447776,0.00413225029818887,-0.0189464147022746,0.0152960402921751,-0.00597174427432889
"536",-0.0107554623157183,0,-0.0140485491193485,-0.00942152963440124,-0.017001015695003,-0.00555286559269386,-0.0385332968911943,-0.0254360015649289,-0.0117635636461226,0.0245768480119914
"537",-0.0097208726116369,-0.0124446482848205,-0.0129534301456042,-0.0253622244948566,0.0097161074885237,0.00284397585000673,0.0642024346979528,0,0.0211966802087298,-0.0111942597399849
"538",-0.0357792715025458,-0.0402440262627926,-0.0419947753809371,-0.0246282637695402,0.00923836894512764,0.000946406709411818,-0.0760513898133381,-0.0362490681416204,-0.0007157463993126,-0.00970331719433548
"539",0.0379103927284354,0.0427784520432497,0.0410960916220613,0.0547882152490462,-0.00104851389373972,-0.00377874107228748,0.0823112768122176,0.027582353870901,-0.0306968168209306,0.0190527660614423
"540",-0.0078728278087703,-0.0288384452566705,-0.0263159132333515,-0.0171636522628028,-0.0115494987523489,-0.00906016919419739,-0.0252287702018757,-0.0278183129569433,-0.0166789923990607,0.0117521957846016
"541",-0.0162617065946635,-0.000836131914668914,-0.0121621122306897,-0.00873157875891872,-0.0105258505106456,-0.0025521779103862,-0.0423854729100496,0.011546503874154,-0.000966226495625944,0.0211193055324381
"542",-0.0223481124746896,-0.00711606344545523,0.00820785947884461,-0.0157628558831904,-0.0057571087721483,-0.000852212882174852,-0.0152760976323317,0.014391907672731,-0.0046206856785016,-0.0118925004637856
"543",-0.0450425156533952,-0.0619731621757258,-0.0352778894428293,-0.0607629919745299,0.0165548825634956,0.0100324948378487,-0.0700081983859879,-0.0631116951787594,-0.0183525537629025,-0.0502355994577631
"544",-0.00750716896562464,-0.00898868813990406,-0.00281317861535169,0.0140425446908465,-0.0066806290408068,-0.00127062639060282,0.0038495036362316,0.00574417938402938,-0.0097877378203014,0.00661170746738571
"545",0.0236906372858814,0.0380953292982193,0.026798407196351,0.0702273879670319,-0.00458130339754625,-0.00508961086410264,0.0264171684155863,0.0150569581317637,-0.0116615169739948,0.0350300751350248
"546",-0.0408474796404067,-0.0397553826765709,-0.0192309336704583,-0.0411274412819459,0.0278108049079433,0.0117233879425833,-0.0643421337646198,-0.0424550464465263,0.033711653752369,-0.00846112494133433
"547",0.00174379512811207,-0.00136511510570436,-0.00280110911372899,0.0168673164164961,-0.0066692535107753,-0.00474013976289434,-0.014640836792663,-0.0186966118757187,0.00326125672923716,0.0240000562089202
"548",-0.0117526884405131,-0.0241456763104482,-0.0351122170728579,-0.0194313211767954,-0.005851041442547,0.000423245424358898,0.0211617001168976,-0.0446379480431427,-0.0186369160403412,-0.00572919525600046
"549",0.0596094133178195,0.0732958877478145,0.0509461451735032,0.0811987469976443,-0.0191992487741059,-0.00730017081536793,0.132275333548172,0.0717948410799516,-0.0268300872253504,-0.00261919038814651
"550",0.00651278667223765,0.00521984670507147,0.00415506591646309,0,0.0108202586357005,0.00714049992520271,-0.0171343273768156,0.0159490316473783,0.012253256322365,-0.0315125524628562
"551",0.039371968675505,0.0359151187798117,-0.00137934570413001,0.0384442983713824,0.00476880120676038,0.00285703913626301,0.0788429855278885,0.0387229781787357,0.0210714747694298,0.0466376618266351
"552",0.00781429999984118,0.00167069034310696,0.00966855079029361,0.00559621715714553,-0.00503633726120079,-0.000739012105462344,-0.0212998834020881,0.0292192167753065,0.00219544461460908,-0.00880838321565069
"553",-0.0030222970778232,0.0104253980193358,0.0177840282909425,0.000855917712214715,-0.0157700043386888,-0.00570179661656423,-0.0735459276597641,0.0234949083488347,-0.00547645107963468,0.0219551233768189
"554",0.0305823454179757,0.0222865850372336,0.0349458852986433,0.0218135584711687,-0.00543893155571729,-0.00191074420633464,0.0745243329816703,0.0325203237692255,-0.00837006580275113,0.0214833462568833
"555",0.0223844930479018,0.0270487056843443,0.0233766849657724,0.0209291058666849,0.0378874897947294,0.0342616848671105,0.0516394592634593,0.031033027465418,0.0338737779445382,0.0125188655265474
"556",-0.0123862799178847,0.00353786180518112,-0.00507612160209581,-0.00655982134080479,0.0012457253681859,-0.00339462788651601,-0.0569893827498497,-0.00628959943268437,0.0135353104967368,0.0207713816451687
"557",-0.0212939139166581,-0.0117508629009405,-0.0216836233156422,-0.0136195381877996,-0.00555079948665904,0,-0.0744964137992823,-0.0134092163216231,-0.0080551353058852,0.0135659568000472
"558",0.0718295707963443,0.0729292343975132,0.0782270795442137,0.0924688277053707,-0.00866032880217582,-0.00340670695439915,0.149897659421945,0.0411020138724347,-0.0161341389522017,0.021032562538039
"559",-0.0197034188389276,-0.0369415577860798,-0.0278115703272275,-0.0310229650682626,0.00951323662710157,-0.00145031391586148,-0.0714285674983561,0.00897250944399919,-0.0122719914797569,-0.0163857844833152
"560",0.0105458251262904,0.0149597767396972,0.0298508457947098,0.0150200948205002,-0.0134623346781926,-0.00601616478857048,0.0138825691193822,-0.00222281786247169,0.0113249701371623,-0.0152308792253397
"561",0.020380732271847,0.0120937187204595,0.0108695194703741,0.0272584211765272,0.0115991056461537,0.00260884886984525,0.0248256930985233,0.016042973898523,-0.000543629032062398,0.0173997215694346
"562",-0.0180489544833161,-0.0403285846846951,-0.0167264053537252,-0.0295677927318129,0.00741847150607677,-0.000624821304657797,-0.040120811304677,-0.00350892812366876,-0.0134885021211791,-0.0185273076455011
"563",-0.0345542459384278,-0.0412452143025946,-0.0388823024085141,-0.0515623778272277,0.00382600739244632,0.00427033146358391,-0.0548108613142988,-0.0528169515972947,-0.0078288563716209,-0.0363020355662409
"564",0.00926511469461477,0.0381491494305963,-0.00126410449317971,0.0218285668709286,0.00714528860492525,0.00176324968054664,0.0621610220656348,0.0250929871978089,0.00333402967323759,0.00452038323437498
"565",0.0193662682770022,0.0234561216670568,0.0291138798100663,0.0330511104246944,0.00912594276203449,0.00245039348960496,-0.00903404961510446,0.0117858060215545,0.00830748790770364,-0.00249996577856626
"566",0.0292374533134969,0.0469822407967126,0.0356706146405892,0.0542334892952243,-0.0122207987667173,-0.00652481164826502,0.0661911621540179,0.0640683531509216,-0.024497374761039,0.0385963742912467
"567",0.00994891974325207,0.00839127941885498,-0.00831360943605863,0.0122129943998104,-0.0204624685571595,-0.0114682355576176,0.0895909322513835,0.00505243830081281,-0.0136262044946103,0.015444053609444
"568",-0.00783316165564696,-0.0188132953445668,-0.021557151427733,-0.0124313912747096,-0.00427564515539114,-0.00232025905529232,-0.0160352357054271,-0.0146626659134874,-0.0264870316925234,-0.0123573436304513
"569",-0.0233256194086409,-0.0265487954133601,-0.00611992672128725,-0.0229545750613867,0.00253774204250967,0.00253718283203819,-0.0752429630508087,-0.0153060769244497,0.0172393696694981,-0.0178056351805647
"570",0.0107778399406058,0.0102273739629903,0.00738946314561528,0.0147783901251968,0.00885652478362453,0.00495524543674497,0.0209975256818271,0.0250429503569414,-0.00149869729072394,0.00734928855250017
"571",0.039742995988193,0.0217475506248983,0.0366745498140268,0.0436894162074914,-0.0125421076852887,-0.0058747237772504,0.119353892353534,0.0421234824712589,-0.00346383785401416,0.0145914913061271
"572",0.000233536288142489,0.0176143823753199,0.0023585512868296,0.00608219609791849,0.00918411373942729,0.00590944010554884,0.0127947605916332,0.00525428790727656,0.0181902333029831,0.00431451718146958
"573",-0.0172438084470581,-0.00937609290186214,-0.00941155091469736,-0.01600282524381,0.00522777739728775,0.00514199839761353,-0.0819564538328632,0.00723736008072406,-0.00580330015259334,-0.0181385200973956
"574",0.0106699983458791,0.0152894945315916,0.00475046720078898,0.0144561821960447,-0.00173342829383505,0.000938762596447429,0.0818630466520858,0.00518970139987673,0.00148789052920151,-0.00631979731497179
"575",0.0146628077738691,0.00609542462108448,0.00354576757420144,0.00854995568322581,-0.00791066246723893,-0.00396289114257808,0.040769613622613,-0.00198528042921309,-0.0193143085714287,-0.00440312116309871
"576",0.00670545924430477,-0.0017821900213203,0.00471172276483567,-0.00706455400821548,-0.010989278776253,-0.00806212596272826,0.0100282574307373,0.000795231090007897,-0.00687562071729675,-0.0073710074952722
"577",-0.041915900182222,-0.0485539519269844,-0.0222744777781957,-0.0487371026005685,0.015142608698713,0.00696654931682961,-0.10704292471858,-0.0588466672440687,0.0203003517918288,-0.0376237562217255
"578",0.0195374750530803,0.022889458873167,0.0119903954268781,0.0213161890920102,-0.00988005095758848,-0.00387863695855928,0.0913825435333215,0.0190115643606736,-0.000690028775964135,0.00360077366973188
"579",-0.0061132856346614,-0.0110051174468814,0.00355466464553267,-0.00842169254219738,-0.00606534642689938,-0.00241943568749059,-0.0337469180217776,-0.00373138862382139,0.00563929112256067,0.00153775748535745
"580",0.00981795227349047,0.031527879309436,0.00590333905164542,0.0155095288937293,-0.000098830820417839,-0.000211189207832252,0.0415154721543121,0.0228880764284043,0.0162509275435201,0.0133059086425964
"581",0.0151105843316124,0.0172602443565735,0.0152581153945908,0.0189092036734326,-0.0100399025678183,-0.00390379146893838,0.0528312928889885,-0.00325467734281892,0.0103603374878263,0.0151515687072972
"582",-0.00946231338865933,-0.0130788639161648,-0.00231240448195202,-0.0335475042586449,0.00427527382624637,0.00413115244474405,-0.0564906102739069,-0.0191836937237235,-0.00791349745972469,-0.0248755890277783
"583",-0.00314550144899128,-0.00286536472722487,-0.0162225539471361,-0.00332354646937882,-0.0163366902697882,-0.00485267097692654,0.0108284123128588,-0.00457707321035905,-0.0141557349925686,-0.00714296929139702
"584",0.0212688332498416,0.0312499111169418,0.00824545344450955,0.0526121525565391,-0.00885687094006904,-0.00540646160609115,0.0396973287843978,0.0292637147710926,0.00660970940170924,0.0231244135623185
"585",0.000343268234756833,0.0045280226289357,-0.00584140945128142,0.00915162871028774,-0.00396129976102311,-0.00170535919508807,0,0.0125914848347746,-0.0120005091814669,0.00351577321474195
"586",0.00537661970996983,0.0124827699287908,0.015276224224001,0.0146494357749045,-0.00688246114384772,-0.00321200920871723,-0.0339391420770027,-0.000401313434282957,-0.0036667813796305,0.0300301367672682
"587",0.0340197648350578,0.0410957307408155,0.0266205024776738,0.0690959964329105,0.00329511837900354,0.000966765360635558,0.0865744878514039,0.0389246638449225,0.0194364814066641,0.0194363296856011
"588",-0.00341094199248282,-0.0108552386407323,-0.0033821056791169,-0.00900324068815683,-0.00123149133403322,-0.000214205082203267,-0.0334872182630492,0.0023176882794167,-0.0043998082626332,-0.014299382269237
"589",0.0173346044933673,0.0216163824367239,0.0237555536567544,0.0171967540770037,-0.00236345446484731,0.000429774729776788,0.0334529130828556,0.0354527370391717,0.0146175750708215,0.0265957801542649
"590",-0.0138916228986453,-0.0179036625557577,-0.0232043221371565,-0.0248805670689352,-0.0244129922362164,-0.0083695993353754,-0.0578038155691539,-0.00744340938448629,-0.00111680811797177,0.00188410047824861
"591",0.0233322866095071,0.0477294759040441,0.0407237051890015,0.0333663143568907,0.00242888732229285,0.00119027816125072,0.0677920236663376,0.0292464512636592,0.00603757812974992,0.024917674809716
"592",-0.0187137279834775,-0.03068640979632,-0.00978240723279322,-0.0234253236595574,0.0142199039792135,0.00940218861535147,-0.0293019563045794,-0.0280512595952243,-0.0032229494368875,-0.0082568156770203
"593",-0.00295911913502755,0.00979110700055186,0.00548825470858527,0.00713150066080015,0.00363445889910419,-0.000642589363487378,-0.0159814470564681,0,0.0112609541473752,0.0101757669694855
"594",-0.025173410036834,-0.0303816672903978,-0.0185590071999955,-0.0366915328363863,0.0108643042385281,0.00460663232393244,-0.0679700039241952,-0.0431030227082859,0.00429987886328154,-0.0114468713857856
"595",0.00857021558011373,0.0103337644779671,0.00111247515418045,0.0143669037776575,0.00389078683692423,0.000107577594725017,0.0319459469629952,0.00940027345270833,-0.000658656302937932,0.00648449018123598
"596",-0.00816156071900942,-0.0131971711200662,0.0100000913401466,-0.00922256306055913,-0.000306052399653201,-0.00245338086250613,-0.0328327753910836,-0.003880357333789,0.00571244650897995,-0.0253106155559778
"597",0.0284072932005732,0.0434636122510601,0.00880087594262102,0.0555184865414908,-0.0155036409907923,-0.00587897405643056,0.0750077368316884,0.0268796951280579,-0.0129983829711071,0.0264399184207804
"598",-0.00120614707954736,0.0124962176578027,-0.00654301534906043,0.0113384733286714,-0.00528422419601726,-0.00139789971076187,-0.015939527519664,0.0170713211454612,0.00664008403452754,0
"599",-0.00669450384299675,0.00474678376000748,0.0131722167142636,0.00311449030678368,0.0105196794025073,0.00312293754643855,-0.0116137236528804,0.010444028264178,0.0141820691972523,0.0160994686754468
"600",-0.0143630170618625,-0.00440950312921207,-0.0130009651833735,-0.0186279111288238,-0.0251492632581566,-0.0109488749408226,0.00185536380626128,-0.0103360779736802,0.0173441517615176,-0.00814846504239086
"601",-0.00212967858099922,0.00379622607312946,0.00329313591519065,0.00442905025506635,-0.0111021527540194,-0.00586083888782862,-0.0212964257291105,0.00522218283558051,0.00319663299300221,0.0146050497443448
"602",0.0256122186970777,0.0211157722642228,0.0328223878122322,0.0119686076938175,-0.0150754220190925,-0.00665891014732556,0.0517183263915939,0.0330236006478395,-0.00414232598741737,0.00224927486095283
"603",-0.0178530435065755,-0.01697528171189,-0.0190676583039537,-0.0115157914262588,-0.0176943316306512,-0.0113205306280054,-0.033282751863283,-0.0114939906935275,-0.00330636725029088,0.0044882691767838
"604",0.0139398275358638,0.0128728032230729,-0.00647951950312986,0.0308563701483406,0.0144773355735592,0.00522422319346827,0.0189204654216342,0.0148979613437157,0.00845372953837553,0.0183200938637791
"605",0.0177080816479152,0.0136391773775599,0.0184783803396797,0.0152720318964594,0.0258167985999238,0.0112798555612725,0.0273970994295858,0.0329399718006802,0.0207979524787341,0.0193066290542936
"606",0.0242084091653041,0.0284403987373192,0.0160085665871632,0.0421177389278784,-0.0295634814059488,-0.0163195214674717,0.0420741838488241,0.0183706919273192,-0.00488559266794986,0.027550648242207
"607",0.000844058853561203,0.00713632513334894,0.00105044705086721,-0.01443421796976,0.00537849362584542,0.00334440092831967,-0.0147852785362761,0.0139554116260816,0.00658098798973183,0.00418930158616559
"608",-0.0126515788363002,-0.0345437204093545,-0.022035646343403,-0.0354419973566668,0.00939112111207874,0.0061122260879376,-0.00230904192414305,-0.0184627618635977,-0.0202365813591056,-0.0333750258162775
"609",0.00939640293952038,0.00795091339598586,0.00751063377411998,0.0185238235093743,-0.0206622742630818,-0.0115963963025945,0.0295054788081492,0.00273566713735773,0.0192776074874437,0.0366854001460537
"610",0.000211691639468103,-0.0127425823865505,-0.011714731630286,0.00208705681927501,-0.00762159953403652,-0.0099459306816978,-0.0126440130428057,-0.0225103028038288,-0.0261873004410069,-0.00541225372086029
"611",-0.00412494800853747,-0.00522438238650458,0.0053880378011899,-0.0154715286863936,-0.00255993313175851,-0.0050791359224962,-0.00369962564256265,-0.000348578981987702,-0.00160069364636317,-0.00251151998290522
"612",0.00509802039540208,0.0120481488208191,0.00857455134963758,0.00181335794803106,-0.000112300070184701,0.00431060557937313,0.00114277869432566,0.0150086467880841,0.00288589146827478,0.00965169779847508
"613",-0.00253623197431108,0.00274722327328325,0.00106253655446698,0.0126696603467873,-0.0157359001848556,-0.00598691936359641,-0.0191156742760221,0.00447043210070874,0.000319716501764544,-0.00374059749461575
"614",0.00444939895516261,0.01674299982856,0.0169852278927056,0.0214476988715422,0.0111124863748817,0.00681879268543706,-0.0186155243620525,0.00581989870843036,-0.00170470912311205,0.00917814283389506
"615",0.00274206909814168,-0.00508986180252002,-0.0010440235960526,-0.0160396438540866,0.00897134795559462,0.00530483416774441,0.0281562814824341,0.00646691218013418,-0.0163286984950489,-0.0140553730163712
"616",-0.0229279352158248,-0.0373158020197218,-0.0177637445657457,-0.0358624668998199,0.00900274491288999,0.00448994562502669,-0.0449694657164911,-0.0246869672122422,-0.0116089836521425,-0.0192872499722414
"617",-0.0135632892237509,-0.0128162949378046,-0.0106386036084579,-0.0150631072587546,0.0174052092868417,0.00558928452742258,-0.0141864998018745,-0.0149100189016231,0.00911088933284065,-0.00384783372232922
"618",-0.00098205858364242,0.0031662917716444,0.0118284254746104,-0.0112358856509557,-0.00563038418245942,-0.00266749085154794,-0.0140841938603031,0.00457605064521882,0.00456867181551179,0.00300442766130105
"619",0.00731850856240679,-0.00315629801122252,-0.00850165348527121,-0.00284084191850309,-0.0151355648036768,-0.0121482197244771,0.00496870996683341,-0.00455520579281143,-0.00801296173281996,0.00128359132876055
"620",0.00368553803250138,0.0145657867521098,0.0160770084384925,0.00506474301412507,0.0137104607043168,0.00462585465606091,0.010815582611222,0.00997173902342308,0.00316560415712686,-0.0085468920092806
"621",-0.0299868946405457,-0.0362211551102113,-0.0221519367148924,-0.0362204562871901,0.00970580442855318,0.0053899857830999,-0.0510548174922851,-0.0278563478586329,-0.0147987047921936,-0.033620804004005
"622",0.000784118507420439,0.0201985666026792,0.00650774566384849,0.00649001903319735,0.0117734072442681,0.00323956133302539,0.00869876466348374,0.00652896244471579,0.00419700680144675,0.017395175235059
"623",0.00861831087304221,0.00194736672680018,0.00215499945380415,0.0219314007476987,-0.0100348940594503,-0.00378539197209382,0.016437945745458,0.00504474140738553,0.00582928961349061,-0.000438398234711701
"624",0.021748184143084,0.0129576231729216,0.023655930830268,0.0297887778793828,0.0183327341404746,0.0125169755876151,0.0159490269705911,0.0340626563199051,0.00940405717017123,0.0087719456635289
"625",-0.00260641324326283,-0.00319775049099835,0.00315152154104514,0.00528769472818924,0.00169419133529969,0.00132457608472158,0.00879123214254762,0.00970852597093641,-0.000216628755641324,-0.00826089106396555
"626",0.00936418279477635,0.0112286631818617,-0.00523563116541537,0.00742584477389086,0.00148066233067667,0.00209423064042746,0.0024895878372635,0.00583823767814051,-0.00270885250071673,0.00964489652745826
"627",-0.00809056634310457,-0.00444187661495998,-0.00736840605180156,-0.0101352974459106,-0.00168948971702554,-0.00264011878996451,0.00651968739341235,-0.0191191611942768,-0.00934377434437439,-0.0178027572355389
"628",0.00413290431183344,0.0152965593370658,0.0116648887971855,0.0183057889121763,-0.00198407634705167,-0.000641125693905065,0.00987055799939407,0.0156629976478182,0.0132704430796227,-0.00397881616864659
"629",-0.0272938486894216,-0.0310735590804828,-0.0220124094871148,-0.0274221657446063,0.00233906792563121,0.00331914381058418,-0.0455098852854101,-0.0215905468403288,-0.0123389870368978,-0.0221926019969989
"630",-0.000111098794276399,-0.00161957086279385,0.00643069971056254,-0.00219275487817117,-0.00190868178385784,0.000661926338197283,0.0208000957498877,0.0091072254651321,-0.00536984109589045,-0.0299592023076115
"631",-0.0193763838914983,-0.0295262188725663,-0.0106496550486995,-0.0235482738638931,0.00669383515883193,0.00396928021781107,-0.0369904839751437,-0.0357513731943744,-0.000550936523778467,-0.0159100812892855
"632",-0.000681352849270178,-0.00668689239904308,0,-0.0115753451365109,0.0184691831682438,0.0115280963990267,-0.00976602840625007,-0.0104394370780957,-0.0158747879602555,-0.0123634141565601
"633",0.00193184402894708,0.0151465299264681,0,0.0178918143645745,-0.0119174556504457,-0.00586168650502361,-0.0161077720259837,0.00800308065981814,0.00268852927148622,0.00625904125719567
"634",-0.00238185769227295,-0.0079578382104889,-0.0107642272585805,-0.0118247561630231,0.00922957663432444,0.00622358791972233,-0.00167067557726697,0.00360858844048839,0.000782035509282908,-0.00765554569948457
"635",0.0243294951656052,0.0257354245007075,0.00217636158954382,0.00711534484047971,-0.00561206787056134,-0.00358078768278358,0.0394911931642492,0.00898948347393858,0.00680955555236551,0.00530393685595221
"636",0.00566023298011653,0.00260693673246815,0,0.0109182326377255,-0.0166161407569911,-0.00664292789644993,0.0115906687079375,0.0242336091474362,0.00687433181340857,0
"637",0.0292464309154865,0.0425737946362419,0.0108576941507599,0.0536848967162606,-0.0257173193517866,-0.0129356694001683,0.0343731680506618,0.0208770742977682,0.0157471647560217,0.0263786816745606
"638",-0.00160840439219612,0.0109101041048647,-0.00429661927371194,0.00180880414289875,0.0107994749074471,0.00599744004854763,0.0129232025740091,0.0248808029248819,-0.00281867959277282,0.00233656119252856
"639",0.0109544117882654,-0.00370017730033678,0,0.0102318322665111,-0.015431827226783,-0.00673460016712224,-0.0233901858288824,-0.00897910479287389,-0.000543629032062398,0.014918402839005
"640",0.0106237128967508,0.0194985607416231,0.0129451280908695,0.0357464719013676,0.00526120886936732,0.00366785173038053,0.0323482955772509,0.0218121531273721,0.0146850756010006,0.0165364813130622
"641",0.0046256465592347,0.00455383732603187,0.00851980606543523,-0.0028763047449345,0.0199520583892705,0.0111848087907211,-0.00210929839801899,-0.0042690964210812,-0.00160808320763384,-0.00361499950632049
"642",-0.000209489844783861,0.00392852443117997,0.0116154290456298,-0.00230757387684022,-0.00897971269048048,-0.00591349781208339,0.000906126301100318,-0.00428757667286983,0.00332873413493195,0.00544224272584604
"643",0.0220825990602811,0.01745963868509,0.00417537044449379,0.0283317150367384,-0.0183363157097958,-0.00969500129836665,0.0346906804077367,0.0215300772688221,-0.00192636982178152,0.0207486147016711
"644",0.00409597672250261,0.00739624063692479,0.00519750382104189,-0.00477908294870544,0.0048347992616169,0.00211363122916919,0.0087461573671368,0.000648759422275269,0.00160842801611771,0.000883861571832734
"645",0.00295720548761969,0.00146843546066133,-0.00206827016296107,0.00875702076182061,-0.0114822355963174,-0.00466217625359167,0.0187865199309125,-0.0116656368032546,0.00321159391021975,0.00397354664689109
"646",-0.00467721802513221,-0.00586500975144277,-0.00103601744676962,-0.00448042575961749,0.00884982454189154,0.00200719015984818,-0.00397172566528536,0.00557366940134196,-0.0170739303924227,-0.0109938289580486
"647",-0.00245171615025896,-0.0097346287188681,0.00726130268981029,-0.0225034758653664,0.00548189296107404,0.000668292242900881,-0.0142411400284501,-0.00912941840442005,-0.00987953523092455,-0.0257892071251772
"648",0.0104455070398519,0.0196604846461275,0.0113284252389072,0.0247480309442458,0.0141772938986904,0.00400441054965039,0.0349609591765705,0.0164526737396815,0.00460532909885947,0.0310360066831867
"649",0.00141879427245462,0.0169441898036939,0.00509164821993391,0.00477385344369718,0.0194621873884144,0.0100817323237641,0.000837576636459669,0.0213660709504782,0.018882284908897,0.0199203653748934
"650",0.0164960879231288,0.0264293138593281,0.0172239238866898,0.0374508745520838,-0.0151548681350057,-0.0106267037208979,0.0198047745467906,0.0288431336120107,0.00557048753230815,0.0282116866853799
"651",0.00258880433823783,-0.003358734691292,-0.000996009735260595,-0.00915925261617978,-0.00795123727622093,-0.00289086288527318,0.0475929516185372,0.00462123557124028,0.0086289227028149,0.00042220018779604
"652",-0.00287956842164572,0.000842532528478213,-0.00697884210457611,-0.00842845488529287,-0.0149484030101901,-0.00568665050854533,0.0404699896240335,0.00275955908250247,0.0010561787072243,0.010548596042903
"653",-0.00517879685459333,-0.00841766083682871,-0.00100400958407387,-0.00822584043290242,0.00340894514452095,0,-0.00627342113600182,0.0015292339328179,-0.00189914540936009,-0.0229646233327346
"654",0.013114087231656,0.000283105201185574,-0.00402010430268906,0.0099529480201539,-0.00832908463635273,-0.00661656968605173,0.0464646555507706,0.00091575716579162,-0.0089851798939784,-0.004700702637916
"655",-0.00207462126147018,-0.00735488546477925,0,-0.01122379436378,0.0124875633130188,0.00643474339921202,-0.0197879186631147,-0.00274508526800432,-0.00874666666666657,-0.000429451290466343
"656",-0.0124768675406385,-0.0108292972653599,0,-0.0188261747615885,0.0115698746848376,0.00695457061863669,-0.0295417998867507,-0.0171307379996957,-0.00150649951576454,-0.0150343792638081
"657",0.0107290307623957,0.0146931426990529,0.00504540599344505,0.00902964729462052,-0.0106823709442607,-0.00278483668988883,0.00659535867385741,0.0289448411458124,0.00172428061510632,0.00523324715238638
"658",0.0076391493826069,0.0167518194310319,0.00903614574295442,0.0173374809428881,0.0141783186035394,0.00781971360040901,0.00478873747297692,0.00574705183213009,0.00828406696990003,0.013449063960312
"659",-0.00767956785038904,-0.00949457411986543,0.00397966113425685,-0.0181414847625702,0.00387166444604214,0.00310356841789661,-0.00902968209105659,0.00330839497561519,-0.00768246897479219,-0.0282533912361369
"660",-0.0246056822418017,-0.0352411298298992,-0.0277499633074083,-0.0391937958847243,0.0147828161054713,0.00685071440117757,-0.0501137337440309,-0.0344723875649234,-0.0149462258064517,-0.0149779951796416
"661",0.00793403884478372,0.018702495166786,0.00815495286177526,0.0218531895441556,-0.00580575677305883,-0.00351190616144126,0.01225715994958,0.0229740161434171,0.00491209469586185,0.0196779575566206
"662",0.00877984954229682,0.00975343707363829,0.0030332580048551,0.00256610531614521,0.00828203375615222,0.00374454558743476,-0.00737069098215914,-0.0145674135376276,0.0051053770390046,0.00701749333334312
"663",0.0103044928347111,0.00909072557790225,0.0120967886434278,0.0173494001790182,0.00821379037905401,0.00263345564305051,0.0405727296142149,0.016322881078056,-0.00280992113703582,-0.00827519375240693
"664",0.0196055915984306,0.0295609091486313,0.0109564316555593,0.0150965792376236,-0.0205764959109888,-0.0101775334276881,0.0221712891020085,0.0148485129270524,0.0149561617521241,0.00746599767470402
"665",-0.0000971754616071463,-0.00136720994323969,-0.00197057651438914,0.0044062517205905,0.0181290514390613,0.00619114458624659,-0.0057342414929602,0.0050760502511249,-0.0139883179073504,0.00174365530253318
"666",0.00194252374436354,0.0076669099696951,0.00789725528947249,-0.00219337574632006,0.00565668102938299,0.00263721791842131,0.0110332735874616,0.00950642120510925,0.00454847323146956,-0.0143603410888363
"667",0.0000970802083810618,-0.0040758473325867,0.000979425791174604,-0.00302315284169741,0.00458245088848819,0.00131487746346304,0.00446417643172659,0.00176627067135038,0.000323404477718725,-0.00264897051125457
"668",0.00222953068111287,0.00818550054663914,0.00293554729711554,-0.00192930637062549,-0.00393953138318626,-0.00273584963604745,0.00790128225472198,0.00793173510376,0.00431082008502193,0.00841077740029217
"669",-0.000193626161351323,-0.000812198367161066,-0.000975748032788659,-0.00524713495745999,0.00458021179344592,0.00230457137756401,0.00661451589486162,-0.000583302344961845,0.00729693084457694,-0.00219496822668053
"670",-0.00889937446530509,-0.00622963414666899,-0.00195311279521482,-0.019711247162584,0.000932268029826266,0.00295646061856547,-0.0124118056927658,-0.00670730298679412,-0.0050069349630254,-0.0272766279455596
"671",-0.0220573156455687,-0.0283454486624086,-0.0146772437155004,-0.0189748768219653,-0.00242027719079185,0.00259444068924841,-0.0510104350997626,-0.0284790234599377,0.0053533189431838,-0.0153776794646028
"672",-0.00379242300011196,-0.00364668692197334,0.00297915716702213,0.0106815181779178,0.0145752738214084,0.00545991001620849,-0.0197353628364534,0.00604424557008487,0.0243876459129362,0.00229675452761691
"673",0.00831514258127863,0.00760150887277455,-0.00297030815220234,0.0199941264099499,-0.00615764289861387,-0.00358417831684432,0.0177483455581839,0.0156203335380221,0.0132030041957998,-0.00504131910971206
"674",0.0140087636290822,0.0192792294989355,-0.00198576156505115,0.0193223819237547,-0.0170338917648156,-0.00599385881899739,0.0119731091413728,0.0201123458233132,0.000718243389270068,-0.0041454986395717
"675",0.00862192158830499,0.0249449342365327,0.00895525450126033,0.0206044365379321,-0.00703711251416339,-0.00230316465290914,0.0321501247193898,0.017106623154912,-0.00102531529811656,0.0185013728514223
"676",0.0076751229999954,0.0117680663830251,0.00394465994519355,0.0053836708295063,-0.00116308918402008,0.000879306074480057,0.0201842620467836,0.0188140740710534,-0.00359230216565753,0.00408723115819432
"677",0.0102182871686902,0.0113665033643726,0.011787715029528,0.0131189773079219,0.0184262420925949,0.00746653197027247,0.0141670741561197,0.0125907758202788,0.00638643373740355,0.00542728758512201
"678",-0.000190704668054043,-0.00313627865835875,-0.00097109778975446,0.000528458234429374,0.005510699282683,0.00294316038422404,-0.00313112235745971,-0.00442124023496615,0.0110542685072959,-0.0130453034291789
"679",0.00486785933459855,0.00498171819246385,-0.00388692900968801,-0.00369735225195167,-0.00992768566409874,-0.00586821168577079,0.0287512448128093,0.00471830498355152,-0.00830127564589267,-0.00546948107058731
"680",0.00417933832430539,0.00391315246559887,-0.00780511721331834,0.011929647817122,-0.00511739484585472,-0.0020770430602749,0.0176136424834465,0.00414374349661184,0.00959578409142292,0.0233729683713699
"681",0.0151343816247937,0.0184512481529386,0.00491653627317845,0.0251506955157619,0.0017841044177056,-0.000766762426252399,0.039003405173905,0.0198073685238918,0.0102123557085469,0.0129871590421937
"682",-0.0014907516832835,-0.00076560185929897,-0.00978476150855834,-0.00536693096044405,0.0125757561385751,0.00493307011135125,-0.00488684270597428,-0.0121392871250584,-0.00570521446480976,0.000441898573175337
"683",0.000637477261368868,0.000766188454604411,0.00494062211067314,0.00282634577453944,-0.00890090147851141,-0.00534555540701409,-0.000223162830878865,0.0060722788446308,-0.00674449392971577,-0.00883775159514855
"684",-0.00252965581876807,-0.00918587027063011,-0.00983286864343946,-0.00871121762823956,0.00229817056295989,-0.000657984462227645,-0.0158517096610581,-0.0148147252938301,-0.00314175540978534,-0.0218456740229847
"685",0.00582408488883202,0.0113310523457915,0.0129098771787894,0.0152495617114261,0.0020832941002551,0.00263465287759823,0.0309229860786864,0.0158729431480109,0.0133183914872064,0.0164083024803074
"686",-0.00831235561240995,-0.00789405509712859,-0.0107846517383481,-0.0150205055845773,0.00301542965984503,0.00218787778434826,-0.0335257035652425,-0.0175439957770068,-0.00842777181554688,-0.022421542462665
"687",-0.01101903562795,-0.0202770018187692,0.000991191752180764,-0.0196434787275049,0.0029024300762599,0.00273113098502553,-0.0330805102583555,-0.0181358311597792,-0.0129515225548613,-0.0128440036923365
"688",-0.00533270305829869,-0.00445378640006766,-0.00792068486179986,0.00421855260339865,0.0127134830542515,0.00403012270844738,-0.000712773819748547,-0.000852584993056293,-0.00563816487017432,-0.00789966405563647
"689",0.0179030528470971,0.0142102108393836,0.00798392299984241,0.0128643359871616,0.00877671079130082,0.00173537573171489,0.0389917825298527,0.0145051051575971,0.000515494845360953,0.00889941747812428
"690",-0.00300971638640612,-0.00155657065293757,-0.020791893087561,0.002332480574605,-0.000910633761974644,-0.000432181228158801,-0.0167050015666546,-0.00616760979937503,0.00391547643744028,-0.00371406505878014
"691",-0.00386788728416798,0.0015589973424488,0.0050555198690907,0.00620677000005365,-0.00091125795858582,0.000758153116122262,-0.00698142642047961,-0.00310306740059008,0.0145745458277737,0.0279589470361863
"692",-0.0248130696274803,-0.0298389535445709,-0.0251505997569924,-0.0272425740361095,0.0136956742607806,0.00752250228185125,-0.0424186248615954,-0.0200906014635422,-0.00971167445041321,-0.00634633504819593
"693",-0.00466134334568846,-0.0090934695047592,-0.0134162634793791,0.000264159318631219,-0.00692069696371767,-0.000431090087061103,-0.00978955948332405,0.00664167661912618,0.00490350398307782,-0.0100365005487431
"694",0.0149283544922363,0.0145750190693832,0.0083684591103419,0.023243884851571,0.000101170950065788,-0.00010771738129689,0.0269404148944312,0.00114759219040494,0.014740235394727,0.0322580997056205
"695",0.0143242053172061,0.0188882916403061,0.0114105614416868,0.0165203918460199,-0.00989721738463811,-0.00323448487488431,0.000240679110203867,0.0157592900981927,0.0246443498296935,-0.0120535907304756
"696",0.00274840461787651,-0.00261133209011211,0.00923101585352404,-0.00101602599426254,0.0117298642416612,0.00638199162610009,-0.00312832334137114,0.0146685559213617,0.000782186163298615,0.00180756951475836
"697",0.00765592131073634,0.0172777671948625,0.0111788800846626,0.0122014906953221,-0.0104849151552935,-0.00365427252088379,0.0188269608877365,0.00917398433979177,0.0125048650595461,0.0198466927695415
"698",0.00609690837097521,-0.00643327403292349,0,0.000752991019056015,-0.0229243058931972,-0.00960028882052488,0.00971365622876386,-0.0024792511181021,-0.00771905642337956,0.00398048486315061
"699",0.00391573232035403,0.00880577961144224,0.00200982885356793,0.00828147060005624,0.00156437026818446,0.0029412124257755,-0.00164245699914622,0.00386665412665965,0.00700118658114302,0.0202642210679891
"700",-0.00204319866320668,0.0023108187218035,-0.00501507326917994,0.00174219567369316,0.0052054805886268,0.00228100569537548,-0.0150412472149393,-0.00687751141080817,0.00675940530628449,0.0112263661355538
"701",0.0172159756875219,0.0217723237007295,0.0110887303889129,0.0322977200781325,-0.0148104218991028,-0.0068270350982097,0.0367454719577496,0.0340716825801475,-0.000767331656103321,0.00768576514257147
"702",0.00365940015548327,0.00777135947957297,-0.00498504333414773,-0.00553534903709207,-0.00462605638345859,-0.00327221918274057,-0.00759486505366369,-0.0048217825676713,-0.0126703685928202,0.0101693954337263
"703",-0.007474601991726,-0.0121888881051806,-0.0180359893991748,-0.0137947722452734,0.00813224975618421,0.00459745336595763,-0.02713393062444,-0.0156123343184199,0.00311101494156141,0.00251683053248986
"704",0.00826530914653478,0.0151095431787405,0.0163266692943511,0.019141240332518,0.00785794971093323,0.00152462214437699,0.0231229596148343,0.0210553559230857,0.0101764198488079,0.0142258758004092
"705",-0.00528279420542133,-0.00297725216753553,-0.00301226669737742,-0.0132436317111891,0.00540518029815407,0.00228456617785944,-0.0186390853587104,0.00107127821196085,-0.00777132281191617,-0.00618816184932824
"706",-0.0089734444777555,-0.00273682980731138,-0.0030210397000684,-0.0053685093597583,-0.00599622072201222,-0.00227935883176522,-0.00783489228712608,-0.00642031753916739,0.00319089157205354,0.0211707498222049
"707",0.0101637140908162,0.00998022158857981,0.00202006951088252,0.00834169645963723,-0.00488911409927451,-0.00293674853853754,0.0224932047846427,0.0123851568081708,0.00163853493975918,0.00812996973268176
"708",-0.0114335211818242,-0.0170455771646074,-0.0231851606753357,-0.00827268820571991,-0.00752535924207576,-0.00491006703619423,-0.0109989198276351,-0.024999711812511,-0.00413779838602391,-0.00362906586020384
"709",-0.0108251675061144,-0.0160845303589339,-0.00309623012421556,-0.0125119197793441,-0.0129541129128188,-0.00570023442751033,-0.00615241831863633,-0.0155482095934538,-0.0157502853560786,-0.0182111281800219
"710",-0.00458306245793294,-0.00740717810958913,-0.00414088338497987,-0.0173912557616673,0.013657090393975,0.00860007000184293,-0.0152381443398988,-0.0135775490196078,-0.0000982034154898281,-0.00700753571954482
"711",-0.0188876553820271,-0.0270201215367053,-0.0103951616139117,-0.0457650400046924,0.00473658990607495,0.00306097208713152,-0.0418280832292909,-0.0410108463849707,-0.010996514698017,-0.0257368123829955
"712",0.021453836533067,0.033060041075766,0.0157564563451238,0.0442500956981544,-0.0108948833340201,-0.00479570804597673,0.0431490350886441,0.0330990297524747,0.0194579464074871,0.0311036398292528
"713",-0.0289734006471863,-0.0358422105021725,-0.0124094065317916,-0.0466885455823985,0.0145106341957359,0.00744751899760354,-0.0191097074781813,-0.0221149727788131,-0.00155811663145167,-0.0252065640847321
"714",0.00733896945659995,0.00743482528050565,0.00942421054594011,0.0149055153049056,-0.00442063786029556,-0.00263115884388676,0.00147968711517499,0.0127569823710971,0.0138495856222527,0.0173801378940006
"715",0.00316315114137744,-0.00764362494821891,-0.00103736846629121,0.00157328423189318,-0.00999463347434337,-0.00230811496158467,0.014282001334851,-0.0031491615581466,0.0241462440831046,0.0141666878942486
"716",0.00258004503506215,0.0143422750655298,-0.00207695295902721,0.0185915585521557,-0.00913894914754476,-0.00275421014710353,-0.0179653500697937,0.0103389750852614,0.00601163823043049,-0.000821681464220014
"717",0.0183950410806948,0.0172823647405238,0.00728421823616232,0.0205652587437533,0,0.000220717862782438,0.0207663957225777,0.00682201579050745,-0.00112040151485349,-0.00534540630864588
"718",0.00262048176917196,0.00205909936923998,-0.00619858270368201,-0.00125921694758158,0.000966072548101993,0.0029823032532228,-0.0154999252003921,-0.000564549375918877,0.00420636555786991,-0.0177759529768661
"719",0.0227759265277814,0.0300539828671178,0.0114345022474192,0.0368222685776973,0.00117754802092662,0.000440973112787679,0.0469865457843719,0.0364405252880127,0.00707439262775766,0.0164141340305319
"720",0.000182630012037333,-0.00274303940326082,-0.00719413924722501,-0.00462204763295937,-0.00181926529600918,0.000770097137745118,-0.00493469715395567,-0.0152630177834202,0.00184857192257004,-0.00496887633467813
"721",0.00511017427359106,0.00175038422260387,-0.00103531284679392,0.00855360277475592,0.00418172059423472,0.00285949149993603,0.0184183172018237,0.0102409550357603,0.0111633823338257,0.00665829530987594
"722",-0.0101682191005408,-0.0107339744818069,-0.0165802085732625,-0.0222923300365786,-0.00181466063980129,0.000328837561339501,-0.0118246996211143,-0.0167125393216689,-0.0126824728591692,-0.0148822347476368
"723",0.00541121639456188,0.0126166249993314,0.00948357629684993,0.017100548928064,0.00459863021388496,0.000767686813516688,0.0133738785207242,0.0189469138896963,0.0141391647180407,-0.000839266802493133
"724",0.0145048586935312,0.0174436272587997,0.00939457576937519,0.0250970002103841,0.0117125434076317,0.00536856572652478,0.0226903191364065,0.00929713245211228,0.0172225171719067,0.0289794580824827
"725",0.00116878295355716,-0.00612294206419506,-0.0113754093084381,-0.00356536994449264,0.00536735246252595,0.00217934125636665,-0.0142628208757526,-0.00623116807224711,0.00304581213954513,0.00489801833895021
"726",-0.00062855820777441,0.000739276935530553,-0.0104600316042904,-0.00787185040250526,-0.00586246376056876,-0.0025011433825427,0.0165365384128733,-0.0073610823064123,0.00250066086897682,0.000812252937989699
"727",-0.0130315284813697,-0.017729907423624,-0.0232560724859066,-0.0185142917507549,0.00179060826426136,0.00119903415319378,-0.0198825105492194,-0.0192256608670601,0.000445461024498828,-0.0142044773407461
"728",-0.0035512216625404,-0.0127847958992523,0.0075759356103664,-0.00416467141582033,-0.000210645373270868,-0.0001092290974265,-0.00760762812384219,-0.00588044764287166,0.00569901142389106,-0.00123505925958234
"729",0.0127024828545672,0.0210763573545223,0.0107409754289889,0.0209102893704922,-0.00126132177876848,-0.00141538318635737,0.0113825359278728,0.00957715595644459,0.0119532404470826,0.00453423541191289
"730",0.00153369245144908,0,-0.0127522813059359,-0.0055419869794564,0.00631589163414747,0.00512522829880391,-0.0146993104330445,-0.00809129716250023,0.00384987309607254,-0.0114896742436308
"731",0.00351411835803583,0.012683456597038,0.0172227125925397,0.0116306421360035,0.00460167558992675,0.0033626480749811,0.00396258477800271,0.0075949149133947,0.0164734589957258,0.0240763949254048
"732",-0.0162508878644483,-0.0348723632082344,-0.00846549375390604,-0.0388022500777868,0.00374923330540389,0.00454148513046015,-0.0283257833272874,-0.0304298645271568,-0.0133768218133213,-0.0113497883869876
"733",0.00337685088837802,0.000763562798468342,0.0202773860030345,0.00971815601307213,0.00238568288590879,0.00161390747673695,0.0375151178366095,0.0129570938259982,0.00504085703182455,0.0110701708064096
"734",0.0123704331395131,0.0218658584955829,0.0345189874417955,0.0286279116012986,-0.0111391404475036,-0.00551420589441287,0.012897052504484,0.0264354369072159,0.0150466794798225,0.00729925362220607
"735",-0.000449147207804312,0.00273737068944824,-0.00404425414547505,0.0040786204486214,0.000839244458488375,-0.0020571542752168,0.0147793661373909,0.00138467397206332,0.0153348359686873,-0.00684387248095841
"736",-0.00782040608635592,-0.00719610875508869,0.0142128641795316,-0.00931907692848499,-0.0103847162079861,-0.00466595395542391,-0.00851450666654352,-0.00940269475389055,-0.00402754656821624,-0.000810606791958768
"737",0.00570761470892389,-0.000249891099231458,0,0.0091655206369412,-0.0106001732066625,-0.00741425057091405,0.026892680272163,-0.00111663835600639,-0.0417017449461267,-0.00811360440726594
"738",-0.00153148814288018,-0.0059999383862267,-0.00800778021670656,-0.00860434041937763,0.00128612280438922,0.00274575060065207,-0.0173857825499235,-0.00475135193131981,-0.00562636483516488,-0.00899800029003262
"739",-0.0110968052680512,-0.022384451885612,0.00302701640766601,-0.018562946841339,0.00149744594982359,0.00350590215665703,-0.00604693573140413,-0.0235886862895844,-0.0190964899735082,-0.00990506872576724
"740",0.00374057648179482,-0.00128648472749404,0.00301811965563337,0.00614088718748018,-0.00459404983396117,-0.00196532023242935,-0.00135169182235229,0.0115040470918035,-0.000991446624374337,-0.0125052544077175
"741",0.00563519142787383,0.00154593827397309,-0.00802399243475138,0.00585966856992859,-0.0114840267630369,-0.00339063973521048,-0.00293347601307492,-0.00625549391057778,-0.000180404192724803,-0.00548755975720583
"742",0.00424794585984434,0.00360039837704096,0.00606687545370455,0.00364044536519725,-0.000108504493610329,-0.00493841435985809,0.0144833337217083,-0.00457789044790624,-0.0135354629128316,0.00509348414873867
"743",0.00684011565220621,0.0112762317626263,0.00100501863241287,0.00677175256601892,0.00119449508018787,0,0.0194065419679061,0.0091981420752747,0.00841564215148205,0.00548978970308478
"744",-0.00464809888075335,-0.0114036637998782,-0.00803225513145811,-0.0103290474067261,-0.00444735235617266,-0.00319823966992416,-0.00919066824587578,-0.00882926325389699,-0.000272124460669931,-0.00461984469599885
"745",0.00152655788012335,0.0110227180631797,0.0151820901828867,0.00582511066802516,-0.00119774170631459,0,0.00596299638220943,0.00373543070691906,0.0125215226614783,0.01729955854448
"746",-0.0120158983287775,-0.0268762398686789,-0.013958038636013,-0.0287161412075658,0.0164704758426828,0.00885148056997664,-0.00636615607612279,-0.0160320675791897,-0.0380858513517646,-0.0153464185073455
"747",0.0056575359514548,0.000260716399815619,-0.0020223517252338,0.00273258219633177,-0.00429286950026675,-0.00493495877938832,0.00773284101504834,-0.00212808876946746,0.0149990782559746,0.00421237281712639
"748",0.0101625473182378,0.00763783109209304,-0.00303928469283254,-0.00123837892240031,-0.0177823935386727,-0.0102503784009741,0.0120584724950052,0.00207351363586161,-0.0183570450213046,-0.00964764890606939
"749",0.00359292908519326,0.00833551411023814,0.00799825554569611,0.0100778107474988,-0.00559503888125779,-0.0044550102793548,0.0106155165904913,-0.00443371117407754,-0.00729311848414538,0.00720032777982405
"750",0.00196893308575752,0.0105915094602502,0.00305180825313744,0.0099032295628938,0.000220188177149083,-0.00044735829072684,0.011289455553092,0.014251402097869,0.00357921265101657,0.0176619629297825
"751",0.00473444977204096,0.00255648387632901,0.00709951822549604,0.0100518715819369,-0.0103692922389302,-0.00358055158280934,0.0126419114791172,0.00146374572086461,0.0169873106432479,0.00578508727199134
"752",0.00213358203967551,0.00484425611228545,-0.00402827723722377,0.00339806273985888,-0.00278715404765673,-0.00269541967216935,0.00359699758137078,0.00555372725386971,0.00175343298492603,0.017666362905564
"753",-0.00141942110737503,-0.00126837402613045,0.00404456988603008,-0.00358103759363482,0.0065966570968492,0.00263976501436036,-0.0143369745281637,0.00784927472901975,-0.00994935025473931,-0.00201862644316708
"754",-0.000355476329329196,-0.00152468063938893,-0.0110777476192624,0.00437122252819178,0.0065758418650248,0.00180060721639164,0.00171184659603307,0.00490306359727799,-0.00502466730227336,-0.00121349249101033
"755",-0.00959814773958612,-0.00865119742805986,-0.00814677280124576,0.0033848575967228,-0.00476215365280319,-0.00483001762429036,-0.0194324721004082,0.00143507671170062,0.00355370803329258,-0.0028351171688914
"756",0.0169599113416534,0.0266936992362803,0.0256674617980064,0.0291567302181714,-0.000889548849870025,0.00248338319943886,-0.00239524392866142,0.021496600975468,0.0232038490952167,0.0251827673620635
"757",0.00264685866240533,0.00100022463171712,0.00600600891839354,0.00725800446594493,0.006457964191388,0.0043908150940124,0.00240099489711154,0.0103812675052544,-0.000910801432309705,0.00118857325538912
"758",0.000704021572481617,0.0012487199879283,0.00398006247005456,0.00209191616582083,-0.0133862561554227,-0.00403561138727693,-0.000435403822863889,-0.00527650486174946,0.0164995902415568,0.0178076370356166
"759",0.00422174841413603,-0.00324258248158593,-0.00891945070094546,-0.00579895417318466,0.00168193194356903,0,0.00893218691833408,-0.00669982246887624,-0.00618780367343197,-0.0124417099344923
"760",0.00332757808418305,0.00800774607708243,0.011999768061989,0.0079326185826214,-0.00044784691327493,0.00123895223233261,-0.00669392087794185,0.0053397834916018,0.00496303013896404,-0.000787390854466552
"761",0.00139641574578819,0.00819274230483069,0.00889332836314916,-0.00208331425862884,-0.00548716362808099,0.00067379388194988,0.0047827894745982,0.00419344285280299,0.0132889912914882,-0.00315212641401641
"762",-0.00932619000334434,-0.0137894159758014,0.00685614624482267,-0.0160056966003524,0.0171174875115019,0.00718913297040791,-0.0168761971726817,-0.0105788224005535,-0.0209127163653118,-0.0213438275954736
"763",0.00844599506491939,0.0114855414687436,0.00583626349818367,0.00306481943066061,-0.0116259032730154,-0.00479596933499316,0.0187064960738859,0.00815995477193932,0.00950314977831757,0.000807826564948932
"764",0.00270445934389318,0.00049353307909783,0.0145069065228649,-0.00258528254177159,0.0140026896058012,0.00470700628037202,-0.00345655114984578,-0.000279512587592512,0.00439302488440885,-0.0052461774260445
"765",-0.0112239912515441,-0.0180115917073583,-0.00190639202344189,-0.0115455410711589,0.00618671924732417,0.00446214464643169,-0.00910456742618249,-0.011725114710717,-0.0104436134110829,-0.0113589960663488
"766",0.0124955350940799,0.010553085537429,-0.000955226957606747,0.0202619621270319,-0.00285532803933153,-0.00177723222183979,0.0199078837783251,0.015536861084368,0.00595341867261934,0.00656544367339817
"767",-0.0101685064385247,-0.0256091049171847,-0.0219885040304547,-0.0240653390219069,0.0101299712736618,0.00344868425333678,-0.0102961286889507,-0.025591056465825,-0.0231348194889208,-0.0187525843160991
"768",-0.0192292373186542,-0.0308752948201553,0.00488766874068824,-0.0301651491827765,0.00457778933536357,0.00365888819816873,-0.0283915650737609,-0.0191264468109423,-0.0144115932731488,-0.0124636054323451
"769",-0.0222918223188655,-0.0234332398756725,-0.0107005589623003,-0.0222167748865835,-0.00173592929608113,0.000883383565149609,-0.022975975189976,-0.018917625164304,-0.00186276422102727,-0.010517487817516
"770",0.00512771751548069,0.017524716338303,0.00786651767064472,0.00732146828419844,-0.00456517273364898,-0.00220733857670441,0.00730600989626362,0.0201720224849005,0.00289264725002591,0.00467680669095438
"771",-0.00419043529499918,-0.00370958512896236,-0.0107315618377523,-0.0208021174646518,0.000328213402847499,0.00199076336546167,-0.00861268619845701,-0.013666571704358,0.000744277984435771,-0.0110028558895792
"772",0.0047570699156001,0.00505333073230063,-0.00591750772388244,-0.00255930991795517,-0.00054585018969866,-0.00231821913127572,0.00914507900793304,-0.00353768111953945,-0.00957604145734536,-0.0145486749141351
"773",-0.0114723229641338,-0.0254037503961766,-0.00992057129367541,-0.00692831000319472,-0.000546703333619614,-0.000331865194056036,-0.00951539707667337,-0.00562130037278874,-0.000469313812722416,-0.00347368256874803
"774",-0.0108688902351535,-0.0119467194937515,-0.0140279828912674,-0.0108530775311385,0.00874240747395527,0.00387378786296022,-0.00663329078966401,-0.00684337151135928,-0.00488358363400876,-0.0113289556147773
"775",0.0155511148303888,0.0200604299099711,0.0101623261829851,0.0269071034388702,-0.00907768990601199,-0.00342873982783387,0.0181904157387589,0.0161774684877869,0.0225556721645497,0.0242397840215776
"776",0.0121034024705258,0.0161638260999319,0.0191149402585016,0.00814069925838501,0.00285279998570731,0.00166505218630264,0.0165083175258438,0.0232901276374482,0.00719888338161301,0.0215144674378465
"777",-0.00498269652069461,-0.00954418493789488,-0.00987186472326829,-0.0058038537165821,-0.0115961038481274,-0.00476580757544798,-0.0115681883513016,-0.0149812251165816,-0.00394025485036897,-0.0122155473463933
"778",-0.0308657470072236,-0.0455032754197587,-0.0189429510840941,-0.045177717775055,0.0158272223616871,0.00824052842760525,-0.0373626262047281,-0.0266160480158677,-0.0398343525253271,-0.0332622435452573
"779",0.00206669589227504,-0.0190687707164856,-0.00203268006032953,-0.0111640947781537,0.00217930721137338,0.00320204463880636,0.0187048395066887,0.00120193936605739,0.00297017333610694,-0.0127923788437495
"780",-0.00721900381739182,-0.0111490041287868,-0.00712807864379894,-0.00994619072955283,0.00130410631511868,-0.000880358591808572,-0.0227217457230894,-0.0237092036997868,-0.00611386129155522,0.000446913439102747
"781",0.0125601569216818,0.0361372096244117,0.00615372709546302,0.0325817030878084,-0.00998880194337337,-0.00539883569108146,-0.00305343636678868,0.02305533079177,0.0131680410114567,0.0178651962283896
"782",-0.00195875343765206,-0.00530114778069601,0,-0.00262929923229971,-0.00954219955480162,-0.00276975916417743,0.00070681841859499,-0.00120188703957202,-0.00275117151119741,0.00394900110499585
"783",0.0104666283691268,0.00729300609233108,0.00509680679755409,0.0263641908979255,-0.00542511089144582,-0.00122132021003751,0.00870987674219892,0.00722020941949753,0.0191209469428955,0.0118007183910438
"784",-0.000832216907147854,-0.00863261356588541,-0.00608528432121891,-0.0125866675613472,0.00411913158687338,0.0023350704277918,0.00910170980712977,-0.00627266830787854,-0.000840063497808186,-0.00561547411050289
"785",0.0157344791633942,0.0230339367713766,0.0102043760199531,0.0257545402558237,0.00188426988010737,0.00221942735015324,0.0268268617757665,0.0135263302855153,0.0241031574728778,0.0304082808699191
"786",0.00473859749761263,-0.0010984699388491,0,0.00355091390665807,-0.0113982545475633,-0.00531478044664124,0.0094596141267731,0.00207555934620163,-0.00337532375364014,-0.00505895277612167
"787",0.00589510366544999,0.00494793902956681,0.00201988605115533,0.00379039259428104,-0.00402960399464225,-0.00356180209125401,0.0133866199322843,0.00562275799211953,0.00668194965675051,0.0088981828450192
"788",0.00207372555832586,-0.000547150216263725,-0.0161288823685576,-0.008559782149268,0.00539458314113683,0.000558869468265444,-0.000219890218935093,-0.00971165156807496,-0.00463722482349815,0.00588001847142516
"789",0.000180009085513522,0.00136843988333069,0.0122948455093081,0.00126958127691945,-0.004135932986021,-0.000781339290467642,0.0041838964707468,0.00267496465138417,-0.00365397822550495,-0.00542802922543661
"790",-0.0121445807892993,-0.021044364453649,-0.00404830797403222,-0.0230788310137293,0.0156037453955604,0.00759774910467081,-0.00789469291907841,-0.00859522883560637,-0.0108187494269734,-0.0163728741687471
"791",0.00919771228521049,0.00949236176100743,0.00203244136729341,0.00960535689209152,0.00243067879109171,0.000554669240598438,0.00972624131949784,0.00956649024908529,-0.00491239229689866,0.00810937083926322
"792",-0.00135377900057354,-0.00884997593814207,0.00202819982355273,-0.00822852086455317,0.00562469106276131,0.00365708998556347,0.00503448487220615,-0.00444184660192581,0.00884870520819003,-0.0169348735900949
"793",0.000632762696562539,0.00502267857430394,0.0060728779828314,0.0101115964513554,0.00515355419266328,0.00154559518079478,-0.0023957978348812,0.00832823000366267,0.010340707420196,0.0176571726432413
"794",0.010384356107948,0.00222073788719723,0.0100605352912233,0.0169405601670971,-0.000438091102626381,0.00103939684399301,0.0102620554582298,0.00855481802666369,0,-0.010156572821003
"795",0.00277053292241636,0.0132963968227231,0.0029880051395057,0.0113579192271078,-0.00131340952453374,0.000551857059577943,0.000432456247064783,0.015209075703511,0.0145298090103263,0.0106884025606933
"796",0.000891400999516012,0.0120285887147396,0.00695169841061216,0.00124778082010479,-0.0025215199311478,-0.000993168003270983,-0.00216056060330838,-0.00316908312223163,0.00549450564297893,0.00972926960187404
"797",0.00302759868397628,0.00135080601102855,-0.00986224263689717,-0.00523432036513605,0.00527496961490304,0.00176799929456717,0.00411349675768702,-0.00115608495779962,-0.00716648769595518,-0.00879774891871954
"798",0.0142935341069943,0.0207712515141878,0.00996047526069699,0.0260584601525413,-0.0131191044265131,-0.00474217666122412,0.0228547765107978,0.0205438306076868,-0.000180492643138241,0.0118343758967849
"799",0.000175023511969297,-0.00396424532497763,0.00690301103588853,0.000732784668097564,-0.00520589601275701,-0.00265983663634772,0.0124368119252334,-0.00481990267272536,-0.00839275351308999,-0.00125311570013642
"800",0.00166275305534769,-0.00159163003865337,-0.0039177773146245,0.00561232844428261,0.000222337409667261,0.00255562933570341,0.00333105697976888,-0.00113941817832908,-0.00145609760073084,-0.0108741776279682
"801",0.00445558338809415,0.00425194903093185,-0.00688291066840896,0.00703750822108073,-0.00256046773060248,-0.00166268672763625,0.00539573640883795,-0.0091275315794741,-0.011392635696385,0.00295987758725458
"802",0.00417507678086304,0.00846767893522582,0.00990095527429835,0.0002405887860506,0.00368382463450301,-0.000887904322381394,0.00495357063776103,0.00690860788150038,0.00119846039274951,-0.00252956316850506
"803",0.000086602153810178,0.00472336337267065,0.00980397377413267,-0.00337250883304729,0.00622712486402044,0.00155553906653338,0.00739304316243405,0.000571713275935082,-0.00598527635332002,-0.00591707919774553
"804",0.000259879169039134,-0.0107077904377365,-0.00485422350566778,-0.00725166379920117,-0.00132678872320313,0,-0.00285422827827198,0.00171450810499252,0.00379809181467605,-0.0119047301272583
"805",0.00796618241569758,0.0163672507196191,0.0097559470795805,0.0129047543699248,0.00796841243646451,0.0038824313571173,0.0259664086323907,0.0168283461899619,0.0188261441599655,0.0133390202979642
"806",0.00592723430842179,0.00285744304183155,0.00386489652255761,0.0108176527007284,0.00428195903775408,0.0012155535878291,0.0121558992285267,-0.00112213232104996,-0.00733701073664839,0.00891716287918798
"807",-0.000512468586096992,-0.00699318721859388,-0.00673736658287649,-0.00761001008139306,-0.00327880670716374,-0.00264812567834083,-0.00393741171481699,-0.00224683473580578,0.00684369036750399,-0.00210443502469138
"808",-0.00506198671817848,-0.0112152590656338,-0.00193802308956659,-0.012940768814997,0.000986255628518506,-0.00132815880332982,-0.0084996467577656,-0.0161984945023781,-0.0186695402816581,-0.01223100333295
"809",0.00534628659322456,0.001318880022535,0.00485436602627876,0.0036418868864192,0.00109634812347004,0.00332407449631966,0.0103666274894938,0.00660899954449712,-0.00489470820922344,0
"810",0.00703339951893067,0.0057955067675397,0.00966177326044404,0.00701507820353475,-0.00470659824963671,-0.00209880660902217,-0.00276231338397814,-0.00256946491175336,0.00529002320185601,-0.00426988417232754
"811",-0.00485483432872147,-0.015453061419083,-0.0162678046629511,-0.0148931309743677,-0.0182563172887569,-0.00996161881413549,0.00316582636326235,-0.0151684589577895,-0.0186484213441653,-0.0111492962624892
"812",-0.00162633947878399,0.000531870858254679,-0.00583677757054313,-0.00268227428688317,-0.00638407632058668,-0.00368863269195852,0.00157354052329706,-0.000871953967924499,0.00451548435045668,-0.0056373907344931
"813",-0.000599770681926959,0.00771089579266704,0.0156557480326001,0.00489004707387708,0.00281720156829346,0.00235596815451267,-0.00357977535966048,0.0116347030913453,0.0169507119025165,0.0017444157174622
"814",0.00634750974901865,0.00949846350947969,0.0125238674678441,0.0180047235147143,-0.00382199563933983,-0.00145454632854602,0.00439090072194981,0.021276381502243,0.00147346906615597,0.0226382280421098
"815",0.000681694503631425,-0.00444314396469414,0.00570907535511278,0.00382405962527943,0.00315954977536337,0.00100864455444216,-0.00198709438138489,-0.00281511606283014,-0.00717240459770119,0.0021286238789695
"816",-0.00340694835443756,0.00656334430982186,-0.0122989679906186,0.00285706758457405,0.00686333154693441,0.00235202155186198,-0.00895879603991123,-0.00959910053556212,0.00907655821916675,-0.000849649729898538
"817",0.00683734660936874,0.0164320700112832,0.0153256100522006,0.0261160851349849,-0.00244528545953349,-0.00207354790983594,0.00462032445368377,0.019384074964369,0.0120239103815671,0.0195577740490089
"818",0.00814977096335823,0.00538857674873583,-0.00283012055931375,0.00902338252970147,-0.0166387318295663,-0.00898206393167456,0.0207953924348043,0.00531318663204372,0.00571374014667625,0.0158465370998924
"819",0.00235763540968525,-0.00689110605000043,0.00283815287411326,0.00298104710006952,0.00160077505128897,0.00294574222009936,0.0201768151556299,-0.000556481765926486,0.00126251241106057,-0.000821006858102935
"820",-0.00571240697224207,-0.0110513790365541,0,-0.00868772932427742,0.0127838601280874,0.00621292115129513,-0.0215057584123173,-0.015863614959035,0.0131495903192793,-0.00369756658899045
"821",0.00346383143818141,-0.00051949932262918,0.00094342891457555,0.0034594250940474,0.00045018761720339,-0.00112202045295062,0.000392488974857885,0.00735266285442182,0.00142238423721897,-0.00164954680753537
"822",0.00656754471291054,0.0145605882389443,0.00282745305834364,0.00620561099357175,0.00236685690071714,0.00112328079697921,0.015889001596225,0.0106681861713136,0.00878825550309359,0.00206531912904606
"823",0.0015891574468101,0.00794463764430087,-0.00187973685174114,-0.00799437436875938,0.00528128723761001,0.0026949046211473,-0.00656509921615966,-0.000555564304473344,-0.0055437962473055,-0.000824475860280893
"824",0.000751693822774513,0.000508306057635632,-0.00188316633578989,-0.00207270612176458,0.00324219837831352,0.00190300947729849,0.0227406370091046,0.000555873127740858,-0.00283160777220404,0.00371290560147886
"825",0.011349108829767,0.0142310267852936,0.00471717227028035,0.0147670930014832,-0.00702074912010009,-0.00268213042447529,0.000949829246288392,0.0127779308437062,0.00301709995532695,0.011508480076293
"826",0.00082548453894904,-0.00350765076656656,0.00469472178742358,-0.00545702221329536,0.00112258612570626,0.00168159634995013,-0.0248716858119582,0.000548269598379392,0.00548529598766079,0.00365708345691451
"827",-0.0159123377652938,-0.0213729377627793,-0.0186915215990745,-0.029263670887702,0.00728669908819479,0.00604039335406004,-0.0208330193996297,-0.0216555227259874,-0.0212054901679632,-0.0182186646443475
"828",0.00377023079409233,-0.00385417157812096,-0.00190510723868609,-0.00400389181650895,-0.0024486061209541,-0.00244636309710744,0.00377771719445086,-0.00504365439860122,-0.000809025544930342,-0.0127835421184697
"829",0.00893075802319054,0.008511865875104,-0.0038165347050455,0.0118233141379931,0.0035692063794428,0.000445768126263513,0.0156498436628725,0.00816699005880439,0.0027889968009176,0.00793648541716063
"830",-0.00181994788341133,-0.00818408429080242,0.00383115644658427,-0.00327173910195155,0.00822613702179043,0.0032317601384233,0.0187244025203872,0.00139652460683903,0.00762604528643496,0.0049731226595251
"831",0.00298348607512766,-0.0108302006462316,-0.00858741319550471,0.00422027173815365,-0.00297665433041794,-0.00233193328785264,0.0145510387067254,-0.00223170048642152,-0.00418486339924962,0.00247419288560891
"832",0.00652770760649379,0.00860234775197388,0.00673705575356642,0.00537008119075999,-0.00353824580868045,-0.00278307668685318,0.0130211757157015,0.00698930539627485,0.0120708695304317,0.00658156363703033
"833",-0.00377629313220063,-0.00155042239243597,0.00669216804480621,0,0.00110968670099099,0.000669628900981323,0.00633395308252505,-0.0011105116483151,-0.0038872867941111,-0.00490381329421719
"834",-0.0236507165704358,-0.0445251968288469,-0.0180438918226914,-0.0357642987186685,0.0140777106257646,0.00937069991765371,-0.031654760826789,-0.0330738728691751,0.0166740310421287,-0.0151951590075315
"835",0.00759630474845263,-0.00487681780195393,-0.00386823771795131,0.00842976018437747,-0.00852643975972855,-0.00508428925816995,0.00344098830282191,0.00632345648533517,-0.00279158168345772,0.00333606789495611
"836",0.0123973274108751,0.0185136715417491,0.0116504898647181,0.0164793293259931,0.00419000631226707,0.00166682011595531,0.041341170662623,0.0159955851024345,-0.000262435487051516,0.00789703081839277
"837",-0.0169615461309224,-0.0155039502880563,-0.00287892480919649,-0.0119825599885814,0.0115279858100374,0.00609912022829762,-0.0311012647470793,-0.00590360331778594,0.00945049010719701,0.00783502902155764
"838",0.0129616971919213,0.00705974798501985,0.00288723694727411,0.00546936966620049,-0.00130685559121446,-0.00262094712426175,0.030966412344406,0.0152714846711002,0.00320736821075451,0.00490995854541798
"839",-0.0235147351676819,-0.040172792615417,-0.030710193673815,-0.0458844541926453,0.0179952847734579,0.0067624057227218,-0.0234429569504736,-0.0406686711934567,-0.0074310894124836,-0.0268729322961048
"840",-0.00595630656289192,-0.0269661730644521,-0.000990220522241292,-0.018096332395873,0.00589268027510625,0.00385359486665693,-0.014066017269593,-0.0153892227114042,0.0019151475080923,-0.0225941773588147
"841",-0.033213604463784,-0.0534063745849577,-0.00594648475066284,-0.0408985736986154,0.0308872068839274,0.0109688428716299,-0.0401370728508696,-0.0551459255618608,0.0295421158933744,-0.0196918202787819
"842",-0.0148751515146294,-0.00579460813889987,-0.00897312934889394,0.00526410105838915,-0.0125015527043874,-0.00271237833453397,-0.0168451219702025,0.00530557243381513,-0.00185670523852988,-0.00524014825566066
"843",0.0440411323696559,0.0763806686291064,0.0281690793975469,0.0720088067259339,-0.0207153053294604,-0.00761537100299559,0.0659140178883701,0.0509161430755989,-0.0059186354760794,0.0193151962987981
"844",-0.00284077507338243,-0.00541487246494265,-0.0225048702743458,-0.0180751801445852,-0.00256426124578146,0.00120615471741159,0.0011347146759757,-0.0141800719633901,0.0262822488730119,-0.00172262936785217
"845",0.0139858812137552,0.0163323634119208,0.00900905746054681,0.0124377927983708,-0.00760446239968415,-0.00251884472749386,0.0162452376345106,0.0107880419887971,0.00613291874248567,0.00819678682120339
"846",-0.0124308562457711,-0.0219903888103642,-0.00793631722899968,-0.00933679085234274,0.00658298975115468,0.00274443887925857,-0.0131973001855984,-0.0103764256245054,-0.00691930795849582,-0.00855803888595574
"847",-0.0181050211785316,-0.0302683023752672,-0.00700000660582956,-0.0205852469488547,0.017371027721885,0.00645885411995284,-0.0308908897821965,-0.017076256553233,-0.00157593731877792,-0.0254639689982534
"848",0.00052671677017635,-0.000594243009317763,-0.00201425688343382,-0.00607770205187574,-0.00368849733037446,-0.00217537344633567,-0.00155477936105464,-0.000304684258915278,-0.00839081145491039,-0.0283436440301731
"849",-0.0136024034000837,-0.0190366680980132,-0.0171545693534733,-0.020891418944602,0.0153392597075823,0.00730334852795567,-0.025501430108397,-0.021646522710309,0.00108911694797986,-0.00136734681240436
"850",-0.00569360177735634,0.0042452354245881,0.00718710874425832,-0.00962813961562337,0.00333359675177158,0.000865617525340534,-0.00839024769988739,-0.00218134553280425,-0.0239350660964945,-0.00912836160459607
"851",-0.0377597455146956,-0.0314009313732075,-0.0152903306090388,-0.0496584022719958,0.0210799475209373,0.00973017279339605,-0.0483476469078155,-0.0371642121815644,-0.006773566152111,-0.0207277302351985
"852",0.0145989749953064,0.019950189148588,0.00931669562067139,0.0323471575632721,0.00101706464343931,0.000535754489490392,0.032387509834775,0.0204346833169284,-0.00535216696658036,0.010348075457902
"853",-0.0128310733772029,-0.0259782093997425,-0.0133333413632113,-0.0104443148455609,-0.00345415527353099,0,-0.0200942610913493,-0.017164428082202,0.0140600155002604,-0.000931085981564328
"854",0.00102125050742363,-0.0015687922664519,-0.00623725184803015,-0.0108253649208395,0.00489304213318631,0.00342452719451969,0.0104624219320986,-0.00840875928452556,0.00445057358612022,-0.00792165449983961
"855",-0.00602858547113805,-0.014142120283278,-0.0125523994260697,-0.000547456439640603,-0.00283993272149208,-0.00202624158764797,-0.00393453625509887,-0.00913273122875324,0.00945807762902118,0.0108030940099144
"856",0.0334983476099489,0.0621614750390327,0.0243645090436448,0.0604983506426329,-0.0226883208036515,-0.00951174044601544,0.0542619160700715,0.0513495848605485,0.00185701863883669,0.0292750765132741
"857",-0.0125496097355028,-0.0204083325621176,-0.0165457431973528,-0.0165201900906149,0.00458091478774114,0.0045321148970352,-0.014986970341786,-0.0159673111993729,0.00160076667620235,-0.00857780778638462
"858",-0.0168235235251589,-0.0119483317127077,-0.0031547445613318,-0.0183728243722889,0.0070288705092052,0.00129269017156086,-0.0194194598774725,-0.0104996872335003,0.00866425829401729,-0.0186703822178462
"859",0.02603928680322,0.0310078951893658,0.00527410355352798,0.0350268138059711,-0.00949955320473705,-0.00570139326655572,0.0220497317503274,0.0369772411896936,-0.00108418810493904,0.012065039772875
"860",0.00344399559980868,-0.00210542100897915,-0.00209830838654534,-0.00361699156511697,-0.00729670141638072,-0.00140675074392993,-0.00259678470044178,-0.00279063501380883,-0.015194523419557,0.00550208235748162
"861",-0.035136910813128,-0.0491259611469024,-0.0189275412089821,-0.0355194771858049,0.0268816847362463,0.0138677951511701,-0.0542760647893109,-0.040733404849735,0.0104272889998924,-0.0310077024594181
"862",-0.0124510096559178,-0.00919188790378944,-0.0160775371012098,-0.0155914755113348,0.00766973521489556,0.0040611080093107,-0.0050825085469729,-0.00842800802045507,0.0192968869989614,0.00188232704909397
"863",0.0107121865950974,0.0111964401340843,0.00980397612574513,0.0229381830251052,-0.00497219995501041,-0.00308705006232979,0.0174543282817263,0.0117683965147428,-0.00403323736987793,0.00798490818368358
"864",-0.00534589530695107,-0.00284697569615877,0.001079197993892,-0.00533894241902411,-0.00112198506646533,0.000106905728736617,0.00502059585516457,0.00387728278973465,-0.00363638016528933,0.0046598644724829
"865",0.0292315436531434,0.0491750017891455,0.0172409603913486,0.0348899934726337,-0.0178678746225496,-0.00928673295471383,0.0418402576889729,0.0379784645776302,-0.0131884292167954,0.0166975025710112
"866",0.00485510833300862,0.00332625953101062,-0.00211856236203622,0.00518654209489866,0.012682466023521,0.006357196004104,0.0103896174202192,0.00186054878044528,0.00874170792013351,0.00136868840960847
"867",-0.00154983128223118,0.00693182699723516,0.00636955459556554,0.000258009697426065,-0.00513262221305122,-0.000856853338854435,0.0118643903562321,0.00185720088580732,-0.00341641524178959,0.00273344776777806
"868",0.0227376705162288,0.0359174215421394,0.017932552893561,0.0301778224958333,-0.00412792173712995,-0.0031072266779526,0.0216928695166847,0.0299659022273429,0.0116220737729444,0.0168104514110876
"869",-0.000356787793834634,-0.00953472624082718,0.00414503843687863,0,0.00569940552516757,0.00279467200329631,-0.0072685049645953,-0.00419891497782177,-0.00545496331027306,0.00223419928982249
"870",0.00160761739383952,0.00554250645363163,-0.00206411550078445,-0.00500758596132256,0.00813903743750033,0.00471670328976348,0.00154129843396489,0.000301575083579309,0.0130474526211677,0.000445917171275401
"871",0.00108409316482638,0.00116029864302614,0.0020683848860894,0.00452961779429417,-0.00163505702832123,-0.00202710133957507,-0.00288576443090149,-0.0067132039883615,0.00762920414062007,-0.00178259847966811
"872",-0.0028640338275151,-0.00663017906918228,0.00722394977526997,0.0172847094756481,-0.00286650349462547,-0.00074871270743504,-0.00713888476423585,0.00214015694414171,-0.0198648779636101,-0.00401780231396276
"873",-0.016515788835205,-0.00923719139352008,-0.0122951764024348,-0.0192072068890259,0.0119087263294568,0.00599138885577388,-0.0281770062174901,-0.00762853298741584,0.00880470146029322,-0.00224111676075323
"874",-0.0031030749614136,0.0066164535159694,-0.00428386140741832,0.00257788552937188,0.00679717103844824,0.00372176653652101,0.000599599963135189,0.00491974751380764,-0.0041169206451277,-0.0166218384377776
"875",-0.0165700970236087,-0.0179265481577885,-0.00314776700412955,-0.0176454599024565,-0.00594530297422902,-0.000847852903963053,-0.0205997832756847,-0.0140757319078199,0.00289380743018963,0.00228421090344666
"876",0.00418907307890137,0.00212961180805338,0.00421054156052691,0.0118038583389997,0.00405450078993996,0.00159056402677904,0.0255196745243569,0.0117938820890231,0.0120362651598616,0.0182315253844831
"877",-0.00315189894655943,-0.00394642836892301,-0.011530485726978,-0.00684730036512371,0.00938931356160055,0.0070944424467112,-0.0114387914814874,-0.00797524268059635,-0.0136038283870344,-0.0107431451285394
"878",-0.0308753601928711,-0.0374887067849086,-0.0243903185412713,-0.0406030022892193,0.0109019876802277,0.00431022132246772,-0.0320747908512637,-0.0281386582352194,0.00148650595380317,-0.0276017606022768
"879",-0.00949991438242781,-0.0072830840782897,0,-0.00665414148962507,0.00672816858858005,0.0014654517267978,-0.00985713628550755,-0.0082722890592537,0.00338091044893818,0.00372261089084946
"880",-0.00445650896148586,0.0169060250784767,0.00326092938562783,0.00723459720311048,0.00157672736712855,-0.000440075218249181,-0.00190646998509092,0.0134741719994957,-0.0381327991452992,-0.0152989615223466
"881",-0.00544980121927974,-0.00470516649971142,0.00433352107082263,0.00425655284380433,-0.00797189365776574,-0.00178231092227787,-0.0191000845205181,-0.00158235982976773,0.0123889011244966,-0.00188311652441298
"882",0.00655601889288615,0.0226916083984157,0.0204968228100859,0.0185429888066762,0.00823543716453079,0.00241563413792112,-0.0194720013929066,0.0117310721791835,-0.0167102374328676,0.00283005256186408
"883",0.0314963842591336,0.0354390152915267,0.0190272695602574,0.0221064645724192,-0.0117098581484074,-0.00314336763236456,0.0476608429778249,0.0363519097752865,0.0104712125916879,0.0225775443640059
"884",0.00989506486460745,0.0104166372031849,0.0020746355984862,0.00483491825883386,-0.00637322731477519,-0.00241789905504197,0.0107411849147796,0.000302568558646854,-0.00441691995879756,0.00919974372801868
"885",0.00746543685300338,0.00147276103581295,-0.00621114188999805,0.0121550159360397,-0.00571138569516338,-0.00263344631732376,0.0131274649056508,0.000302425084459212,0.00981146668212163,0.00182312908320581
"886",0.000648567465201477,-0.00264699371596189,-0.00520854904171719,-0.00800604073706124,-0.000403757220391099,0.00168985114737064,0.00370254164154415,0.000906533507590401,-0.00861781844695997,-0.0113739613018505
"887",0.0150882409275654,0.0253612520560453,0.00523582006731149,0.011601236223721,-0.00857041437749639,-0.00495646351872492,0.021926345310453,0.0132850279775063,0.00869273082300093,0.0161067811886209
"888",-0.000091220882607268,0.0025882985444825,0.00729137353099185,-0.00199433399059357,0.0100684642991895,0.00498115241897068,-0.00581496165057582,0.00327776370327237,-0.000506911114338315,-0.00181156937638549
"889",0.000273345352520549,0.0100401331944506,-0.00827279970292638,-0.00474650144283328,0.00996781056592178,0.00516744311516026,-0.00221890300043293,0.00207875662330892,-0.0005917159613259,0.00952804655642714
"890",-0.0275344743989171,-0.0312410883207465,-0.0250263109382226,-0.0298694853229787,0.00488482673198587,0.0057712285322189,-0.0307255070479144,-0.022228721893189,-0.013194662610302,-0.0125843292251807
"891",0.00590673095128125,0.00586352739914209,0.00320873996857629,0.0131956991007267,-0.00615067354868737,-0.00260831398507644,0.01147008059008,0.0142468180093807,-0.00805686994183386,-0.000910226211123244
"892",0.0110914863959788,0.00204003864866631,0.00639630118405954,0.0234932015014728,0.00149745856249539,0.00104586261001027,0.0171137934406322,0.014046851362076,0.00794952887022737,0.00820039019244789
"893",-0.0129979794129115,-0.0171612232159195,-0.0180084068010308,-0.0102296893561314,0.0169436706515633,0.00637354909496946,-0.0192583147540774,-0.0132628262641634,-0.00685815676196899,-0.00271126125667331
"894",0.0223219722030379,0.0361053390073698,0.0183386567927388,0.0302494303623597,-0.0115652071176485,-0.00550262366921661,0.0359650674677281,0.0280765098033497,0.00871819609353808,0.0199366670670988
"895",0.00867898670784939,0.0131393565202409,0.0148309993871276,0.00685092276454657,-0.0106102602816582,-0.00323635572756764,0.0117719372120015,0.0136546739801038,-0.00658912368142117,-0.00310973207646137
"896",0.0104156657960812,0.00733009808816965,0.00104370803522813,0.0068044557174638,-0.00170334820953089,-0.000314026296194592,0.025833465674646,0.00917166414723769,-0.00490997518855973,-0.000891345105075714
"897",-0.0000897432484727734,0.00643727197095423,-0.00521376791936368,-0.00168928461433548,-0.00963747888987032,-0.00345678044639108,-0.00019246907275805,0.00198808137163842,-0.0173995416568441,-0.0107046737841719
"898",-0.00645443185802685,-0.00834293512832751,0.0115303635085287,-0.005560972748342,0.00324314353790012,0.00430970684237142,-0.00153851048338305,-0.00935369704886824,0.00237861858199961,0.00405774690872085
"899",-0.00487221156154205,0.00224356917164492,0.00621757879893137,0.00170196284496682,-0.000302758955530114,0.00209386026883918,-0.0088579203574668,0.00457818051783332,0.0044823519465842,0.0143690478374703
"900",-0.00018138863676187,-0.00167894706013272,-0.00823919939453932,0.00485423840646981,0.0155650610165379,0.00585004868370453,0.00349752310601725,0.00113916998700225,0.0104995799238814,0.0132802587701601
"901",0.0225809824879628,0.0369957360861595,0.0218071667400843,0.0258455454518951,-0.0140379808931571,-0.00309279787466843,0.0303969324731104,0.0301565881897876,0.000432963900475647,0.0192223290506586
"902",-0.0047890651946968,0.00135107236552923,-0.00406529244650511,-0.00470922398077223,0.00577240907981502,0.00470043437619516,-0.00526120372846672,-0.00856122438760465,0.00389472906443888,0.00342901439923127
"903",0.00668314308022633,0.000809791919815783,-0.00204064581456431,0.00141920845710164,-0.00765219746198231,-0.00415810210573875,0.00321106496349155,0.00334268884715105,0.00629367197678543,0.00854337299574337
"904",-0.00106212773180636,-0.000269332519901244,-0.00102248379452896,-0.00448816693291654,0.00466786498234528,0.00480178245823604,-0.0124269979951666,-0.000277645279837091,0.00222757023451359,-0.00465902280095076
"905",-0.00407605468621686,0.000539593520220372,0.00921213106320007,-0.00142402217318394,0.0109057435107751,0.0065454274291139,-0.00324106372076916,-0.000555397049470496,0.0073516240207312,-0.00893604810459558
"906",0.00533875431026498,0.000808562304690064,0.00101415794647508,0.00522813341185557,-0.00369568047298374,-0.000206817537579451,0.00994631900184673,0.00611281030780808,-0.00373382565287939,0.00343490326253937
"907",-0.00539901080885385,-0.00673480388665426,-0.00607922582833265,-0.0137117169304899,0.00210550776018548,0.00505912624512561,-0.0077654028617502,-0.010770874237723,0.00281091136608325,-0.0106975486074448
"908",-0.0274068210731768,-0.0461078766763443,-0.0336391344624051,-0.0318790498483933,0.0134070141010978,0.00564955493832486,-0.0240502764833475,-0.0337795985014503,-0.00331272394514415,-0.0224913537169457
"909",-0.00613047802443645,-0.0025591610839677,-0.00316449176848399,0.00173290271250992,-0.00246766059203629,-0.00255304570194326,-0.0115390898991135,-0.00115597475675688,0.0121868165054311,-0.00752215774694576
"910",-0.0029453432817711,-0.00427581063121185,-0.00105852877239876,0.00543734550125019,0.012471776818193,0.00430044554976194,-0.0021766422604419,0.000867922292070666,-0.00025258062438116,-0.000891650799776267
"911",-0.00046168882521902,0.006011825259151,0.00741579303736439,0.00934144250607916,0.0250268635406961,0.00724001172565591,0.00099158228918883,0.00289010191751893,0.00833758646349314,-0.00312356292659821
"912",0.0122851460897002,0.0108141275230369,0.00525738098908923,0.0104725137357016,-0.00572274643742143,-0.00506135312077494,0.0217907379803199,0.0193083862951136,0.000167017451757623,0.0143241167204717
"913",0.00182508622804733,-0.000844747131048207,0.00627623457270077,-0.000722885644311777,0.00268584756311863,-0.00101779656275025,0.000193917054694737,0.00452347643648943,0.00392485177453028,-0.0039717927589521
"914",-0.0173967375900055,-0.0166243688050208,-0.00207894891135552,-0.00771855290293599,0.0155939139743775,0.00448111243101112,-0.0226788280418829,-0.0115393379948411,0.00141405754937574,-0.0101905157808873
"915",-0.00324424319956895,-0.0160458833102655,-0.00937489638406663,-0.00291667832036757,-0.0011305044404053,-0.00324461476031634,-0.00297513827757234,-0.00740327972083998,-0.00348864526529324,-0.00626679242697858
"916",-0.00381328468011399,0,-0.00630935373299968,-0.00902017901477237,0.000188796946611225,0.0013226603589509,-0.00477406767438537,0.00143442116804349,-0.00158374592328292,-0.00675680343109109
"917",-0.0148428207379685,-0.017181134892331,-0.00105852877239876,-0.0127917022160695,0.0160286517178843,0.00792434201819159,-0.00439757596238188,-0.00888003261827741,0.00484222745735696,-0.0113379006567939
"918",0.00388494606286716,-0.00088897135024868,-0.00317740741390315,-0.0064792588314041,-0.00324801642196237,-0.00453574826132885,0.0130497332409998,0.00780358314223784,0.00830840803997668,0.00504599179799725
"919",-0.00670189019840139,0.000296796213660189,-0.001062811279256,-0.00627040256392808,0.00940312082564754,0.00455641501280102,-0.00554908929675446,-0.00286801912242751,-0.00329599535847069,0.0114102993379197
"920",0.0154898912154586,0.0195670455937351,0.0127659091508847,0.0219587278280229,-0.02831572588427,-0.0114909850315192,0.0159427374846526,0.0192696137007056,0.000413384593364707,0.0171480117157852
"921",-0.0145047595181299,-0.0171561926557878,-0.00315131762499032,-0.0165470909200733,0.0191740882773228,0.00764774678698465,-0.00921937863054612,-0.00846504423662964,-0.000826361444072998,-0.0017746899064317
"922",0,0.0056213285570943,-0.0115912057686592,0.00602687876587704,0.0110835939029412,0.00445265840072429,0.00930516648357838,0.00825281249286247,0.00967660211143473,-0.0133332888102071
"923",0.0299116741194958,0.0385407357049916,0.027718713900601,0.0351971097178938,-0.0206768685679306,-0.00720100031629223,0.0315806930999301,0.0273777919033438,-0.00319462642210622,0.0198197805590823
"924",0.00931201840432738,0.00821529907113039,-0.00311205922951452,0.00168797957587818,-0.0105660821695434,-0.00417122146398363,0.0125502051542983,0.00576935271226198,0.0049305529635868,0.00706713234755285
"925",0.0129713918693422,0.00983397307762957,0.00728378633741444,0.0117956510395381,-0.0123951513997992,-0.00572039186649143,0.0131452405534558,0.0106522998573211,-0.00351623187900707,0.00526322156738601
"926",-0.0112718879560237,-0.0178072152762699,0,-0.0145131691803174,0.0204673054676956,0.00791070901858371,-0.0139013859936201,-0.0132428007520971,0.00689312319962965,0.00523562019718837
"927",0.00702270350649026,0.007365361892818,0.00206639461837632,0.0108642392553024,-0.0079468441927476,-0.00275231645278995,0.000563740720094019,0.00520389668295773,0.0000815158944136307,0.00217010912772109
"928",0.00461928124682465,0.00899884432611797,0.00309271934553856,0.00573200284740794,-0.0197407605693147,-0.00786999698371083,-0.00751428542897503,0.00844687423038604,-0.00937169757453915,-0.00563024417114466
"929",0.00504887750079019,0.00641028753881723,0.00719395601643402,0.00356205483580196,-0.00457259789108211,-0.00288494686813967,0.00397476874637048,0.00162112501896972,0.00139852749915326,0.0104531334813114
"930",0.0111226568737055,0.016062000517312,0.0102045378083124,0.0238997212064158,0.00488667531960552,0.00475329268569546,0.0156488169683597,0.0148370803035309,-0.000903639179241633,0.00732757416011309
"931",-0.000620857250840157,0.00953950231126832,0.00303032819113835,-0.000462193149210033,0.00962821942423298,0.00503860875701401,-0.00297035422874692,0.000531445317460966,0.0197335466271942,0.00299525195401307
"932",0.00381714935328414,0.000539959362641174,-0.00201448718816566,0.00138733382164635,-0.0148343734660331,-0.00347913030449376,0.00781985055563439,0.00106278266692605,-0.000645016948355503,-0.00170654908078371
"933",-0.000265621478462541,-0.00215867185548591,-0.0131179801687248,-0.00507973960883223,-0.00987615401730046,-0.00349157605192818,-0.00535764436075981,-0.0037155165874827,0.00556716950835612,-0.00512813520556832
"934",0.000373624428419816,-0.0102758735525861,-0.0030675407980153,-0.00162440515485995,0.00404893222545399,0.00226754706379673,0.00297232880672182,-0.00583079661030839,-0.000722105449460941,0.00343637901994409
"935",0.0152903256228347,0.0193989280232596,0.0174359484286253,0.0158065413526796,0.00580312867926525,0.00308426992015431,0.0224069713799984,0.0172970841224029,0.00264976712180998,0.00813358273024756
"936",-0.00201374192376091,0.0026802593837294,-0.0110886775977176,-0.00297514222772555,0.0138862700006825,0.00932727273971401,-0.0157578214548371,0.00239155502953081,0.00912948644679701,-0.0106157845556669
"937",-0.00491310411092305,0.000267415330798437,-0.00305813014536649,0.000688797238427741,0.00897021366778006,0.00152197808462495,-0.010305531393014,0,0.00150777713661165,0.00600867863313748
"938",-0.00811161305047836,-0.011758507982219,-0.00408999478773486,-0.00642195338898288,0.00286784030729992,0.00142012234858568,-0.0224324814202916,-0.0108666956468099,0.000792440589360677,0.000853142814789987
"939",0.0206221854719422,0.03163890952696,0.0133472670440409,0.0184672062548359,-0.0134401384532086,-0.00496066966447295,0.0272450428559448,0.0262589594511176,0.00308787799474564,0.0153453669436308
"940",-0.00479018951869747,-0.00655317907483377,0.00506562282775347,-0.00181321026638681,0.0173911030231728,0.00773247570257318,-0.00989903718137641,-0.00626609765880382,0.000236790587468727,-0.00671712532960733
"941",0.00350059323068952,0.00897101811986567,0.00403239064876781,0.00726618264917667,0.00683784317700842,0.00333221598840794,0.00264080421030077,0.0105095128512624,0.00891727423518573,0
"942",-0.00174398614035287,-0.0047072037787419,0.0050202008238367,0.00338138215219974,-0.0041505546377032,-0.0024157255015389,-0.0073378258609228,0.000520150136036124,0.000782158792055565,0.0131023214391592
"943",-0.00297056402657025,-0.00551769917028855,-0.0119880828243185,0.00584136752952835,-0.000663457560098668,-0.00120984478622055,0.00227447613186826,0.000259961999763414,-0.000312567416472787,0.00584064025226727
"944",0.0042060951710603,0.0105681523103975,0.00202198661393216,0.0147418683601708,-0.00483187717732192,0.000535686034651706,0.00491682604124044,0.0161082315354431,0.00781799678467676,0.00207379995796053
"945",-0.00750378167713095,-0.0138563431980826,-0.0191724348168922,-0.00308149840497129,0.00258077172015181,0.0035415164648589,0.00846827274698203,-0.00946077614515217,-0.0034907841597771,-0.00331121313906824
"946",0.0201318676376967,0.0291624239664614,0.0318930467844596,0.0181054265873093,-0.00600678638821017,0.000202241153851368,0.0130619896545134,0.0216832161481562,0.0196948300026172,0.0203488153415423
"947",-0.0000862964021779433,0.00566714026010628,0.0109672985443989,-0.000433752386613806,0.0125657853780146,0.00645157147495978,-0.00294673433400294,0.00757940234014542,0.00625996617070146,0.000406994849060593
"948",-0.00120659341072182,-0.00179297359243713,0.0039446717968501,-0.00889555674455345,-0.00833640024396964,0.00100140323572195,0.00221651700592829,0.000752251531515702,-0.0109248389488635,-0.0101708574073451
"949",0.00560870299651084,0.00487543243043231,0.00491147994297214,0.0120404332777733,-0.00439440398610669,0.000400400499863673,0.00129020880070141,0.0065144418759715,0.00989498388797205,0.0332921999423756
"950",0.00094401000430322,-0.00229840928491554,-0.00195498438386033,-0.000649561821143396,0.000191584451594062,0.00100026750917825,-0.00147229278601058,-0.00174241255870622,0.00478496871380951,-0.00477328649540332
"951",0.00308626478232377,0.000256087249669301,-0.00881490492568404,-0.00411210544642204,-0.00988067268225434,-0.00289811913638705,0.00866474922235283,0.00324200027933053,-0.00249441391987992,0.00479618003680238
"952",0.00777707657470006,0.0174000511435404,0.00296425041358894,0.0184742624928946,-0.00155021348969353,0,0.00987037625653686,0.00870025280002218,0.0159896929984249,0.00477332743478698
"953",-0.00390091390307501,0.006036180565266,0.00689670719924051,-0.00170726652359032,-0.0149444464862504,-0.00571160592688491,-0.00307657099209024,0.00689973235447439,0.00507192484893348,-0.00158359108553852
"954",0.0020430409037111,-0.00249961638537677,-0.00782758905414171,-0.00128238457380958,-0.0122154300564699,-0.00433354667307606,-0.000545073311640332,-0.00587392368527884,-0.0079406827458256,-0.0111022708620921
"955",0.00492782785412693,0.00375944874077772,0.0069031900178087,0.000427984198095199,0.00807833538915514,0.00475738355219324,-0.00508601680798471,0.0078782159863644,0.00448837545944514,0.0100240858846563
"956",-0.0131040491155954,-0.0269664138938888,-0.00881490492568404,-0.0316647719630234,0.00603487668536262,0.00342526108639229,0.00492957298414942,-0.0315093825047001,-0.0310544982950141,-0.0293767432883081
"957",0.00976590427232438,0.0197587111434996,0.00790505181569512,0.0159080206399234,0.00216358618272627,-0.000602608334384303,0.0199854869160263,0.0214372493957653,0.0092998692698496,0.0237218936144195
"958",0.0022054591985452,-0.000503140776916045,-0.0127452168321784,0,-0.0118738234382684,-0.00552554735609534,-0.0019593691553984,-0.00864195666257472,-0.0140877695810663,-0.0123852560833844
"959",0.00186245492739601,0.00075502461905308,0.00794441974505511,0.00108756686278655,0.00675284192185122,0.00030288571372572,0.000178416705830742,0.00498136983299369,0.00200814859034404,0.0084953217711945
"960",0.00295732133068638,0.00327052252051452,0.000985182346324942,0.0108626301737067,0.00286062700124567,-0.000302794001748263,0.00196286561190484,0.00272633801549493,0.00863339269662822,0.00521452919396115
"961",0.000168410639778571,-0.00802404426394199,-0.00984238538390314,-0.000859542681096448,-0.0154416306834898,-0.00666742500238748,-0.00587688435745526,0,0.000229262503816718,0.00518756107376728
"962",-0.00286360437707922,-0.00910017759455184,-0.00298204597787133,-0.0169931590021656,-0.00879130368327818,-0.00579687983324773,-0.0100326527714049,-0.00543742949119286,-0.0103912052876222,-0.00317590168457615
"963",0.000169028599848575,0.0104594023990416,0.00299096517353714,0.00634584909722125,0.00272126960691699,0.00583067958213146,-0.00615254202703253,0.00447308592456741,0.0132798096578193,0.0051772725314605
"964",0.000759874679004735,0.000252529308628846,-0.00397604198699419,0.00282678678649595,0.00934747915965417,0.00447500698438552,0.00072840046301903,-0.000742285754512517,0.010515010266877,-0.00237718728795866
"965",0.00033758082394586,-0.00631010632471185,-0.00998016319365225,0.0110582992357275,-0.00430589899246792,-0.001674731323139,0.00727767184195161,0.00396143253965886,-0.00527821615435886,0.0063542032704953
"966",0.00793056361981037,0.0182879883078753,0.00705652202236839,0.012438042045555,0.0131432394132018,0.00335546223807714,0.00559987975583298,0.0133168384997551,0.00432085361311185,0.0090765567807225
"967",0.00401755845135909,0.00698435139687681,0.00300305776704235,0.00614277444203215,-0.0204000743124513,0.00324132184032844,-0.001077855580635,0.00219021529950325,-0.00694390493833852,0.00469301607448758
"968",0.0192583393100711,0.0240277576284647,0.0229539855270935,0.0227369757956686,0.00778471093848632,0.00807972896592757,0.025894739861348,0.0182125543879808,0.0338982424771019,0.0237446438397573
"969",0.00376229083227431,-0.0128206045153749,0.00878050617176118,-0.00185253040570332,-0.0171530303849617,-0.00420796343209173,0.00999140427712319,-0.00310005893399401,0.00257300597348387,0.00418253064980045
"970",-0.00187432511642849,-0.00833120158548339,0,-0.00412482915765822,0.00449013694761913,0.000301745181287005,-0.00485953515431148,-0.00956959389299095,0.0102653904434158,0.00265047491442716
"971",-0.007184252135363,-0.010377910529408,-0.00676978044298193,-0.0126320539538284,-0.0220477783317533,-0.00844818765401423,-0.036100407623938,-0.0164250051784457,-0.0158949268100952,-0.00679756808052623
"972",0.00402942297856135,0.00124808255082787,0.0116845606292368,0.00734058155227002,0.0013499839415283,0.00375289217427288,0.0119412686175449,0.00171883545822249,0.01216910575025,0.0106463598290467
"973",-0.00376743853440764,-0.00997484760503198,-0.00577486037398656,-0.00978546707123573,-0.000518457496153979,-0.00111176202469243,-0.0080457419612231,-0.0132384888322246,0.00306032486664498,-0.00827682583247247
"974",-0.0118383354092407,-0.00554175374992771,-0.00774446220667913,-0.0241797679262798,-0.00539811149475211,-0.00829522809063132,-0.00937263110828246,-0.013416055359865,-0.0288391826575858,-0.0417299075536764
"975",-0.00141405249466653,-0.00202598450419589,0,-0.000431238585529958,-0.0208746842097293,-0.0128532598156396,-0.0109172294473427,0,-0.00949961837834368,0.00158342810595902
"976",-0.0155796433326655,-0.0253809586058716,-0.0175610976579705,-0.0262990386988423,0.0248371637628892,0.00744062734494544,-0.0314565480031378,-0.0198943926970796,-0.0109499850619239,-0.0296441914335533
"977",0.000508030061691089,0.00364574750559443,0.0148959172811451,0.00509243320727371,-0.00551296039682736,-0.00287159629648837,0.00873665629172082,0.00179894271620373,-0.00450481786283241,-0.00773932753243955
"978",0.0147180774465563,0.0238715205682025,0.0254402633801007,0.0237882775835598,0.00407954048120951,-0.00236679208641832,0.00696668651260302,0.0159013971613831,0.0131154389816137,0.0270935643193935
"979",0.00275105940375253,0.00380133533778726,0.000954188096101705,0.00064556784609171,0.00614583897774423,0.00206228508831829,0.004674341643645,-0.0053018254697883,0.00083277313446195,-0.0143884167031987
"980",-0.000831253164949586,-0.0143904049792994,-0.00285969652977014,-0.00301012732086914,0.004244503918031,0.00535119455953081,0.00204754518939043,-0.00380699327275358,0.00968229220156491,0.00324407562208728
"981",-0.0144769181877274,-0.0330428161620526,-0.0191204429592833,-0.0317015256288428,0.00494861864246499,0.00204717302470203,-0.0070581119665597,-0.0236940978008761,0.00696739607334118,-0.00242518921933998
"982",0.0147737322873818,0.0105959340503494,0.0175436657604213,0.0231622193676602,-0.0178499449990768,-0.0107258305904748,0.0192668569762398,0.0120040872962606,-0.00171126399192723,0.0186385273102563
"983",-0.0116469915236994,-0.0152030765155502,-0.0162834597294108,-0.0248146905786233,0.0138919652060203,0.00433728264889721,-0.00293623035710588,-0.0128933701526621,-0.00797430359084894,0.00477332743478698
"984",0.00303041044190078,-0.0167690197739486,0.00486863788576541,0.00781269425174647,0.00855030515047939,0.00215885363559098,-0.000552206843193237,0.00261235610476174,0.00300498833292018,0.00197938699468603
"985",-0.00562294168534505,-0.0151596843935038,-0.00484504909617733,-0.00819518551117593,0.00520944980238025,0.00174391877283964,-0.00386742708213239,-0.0122459626990582,0.0143060674970439,-0.00948249177806404
"986",0.021267835810679,0.0321605366586462,0.0204478533787145,0.0285843520282469,-0.0222294135375596,-0.0131506809181619,0.00758004225649112,0.0269055024872875,-0.000295325657883816,0.0295174429557872
"987",0.012808497301058,0.022902870610759,0.00954199221713381,0.0197567175372309,-0.00260680211650199,-0.00249647353539573,0.0135778254228274,0.0215774801775179,-0.00132964982531958,0.00852383101731813
"988",0.00269255097707743,0.0119758980969942,0.00567104333923307,0.00361929880235912,-0.00784219353127269,0.000104431408372463,0.00144828502840189,0.00578329826441082,0.0212278850864176,0.0126777038589156
"989",-0.00105768402777084,-0.0100335274974481,0.00469925193099119,-0.00169704811419891,0.0141220975213616,0.0062562446986234,0.000542222223587796,-0.00400001397161598,0.00753236725772033,-0.00113815050425914
"990",0.000570340226719868,0.00571766128673734,-0.0121609296649855,-0.00467475067333123,-0.0214064434448999,-0.0165802134923401,0.00325203093897897,0.000250831153511433,-0.018762137741628,-0.0068363323991949
"991",0.00366366868553225,0.00594290655403618,0.0028408231442123,-0.00640493727427993,-0.00966407172867201,-0.00853533958312891,-0.0149468258017239,0.00250969209677665,-0.0125275238095237,0.00764819747851098
"992",0.00389339426672453,0.00154154036789533,0.00188874652894411,-0.00343782707088336,0.004932652912641,0.00212588237875488,-0.0107858758198394,-0.00150207970588778,0.00430300489740354,-0.00265651027620528
"993",0.00581784072893066,0.00461581034122971,-0.0028275453134603,0.00452795270883555,-0.00608158997240049,-0.00848504299969033,0.0103492369067117,0.0035096695203225,0.000295552939925781,-0.00152208837496137
"994",0.000642682318822585,0.0104678218261363,0.0132325079279085,0.00643909533651832,0.00375665372933986,0.0032099924137039,0.00256061897418047,0.00949289839482148,0.00472637900520279,0.00990851900668721
"995",0.000883083161401066,0.0015158574078884,0.00373157461278462,0.00149278819853871,-0.0145454146443545,-0.0105561069364941,-0.0102171428441464,0.00445405844642521,0.000955457531301773,-0.0026414734242225
"996",-0.00457252289890753,-0.0151362632980371,-0.00650582903361585,-0.0161844034804673,-0.0130229716998966,-0.00409468630257748,-0.011059641325557,-0.0101008574564991,-0.010867940050489,-0.00264846928545504
"997",0.00580205868026762,0.00512297489583391,0.00561298846971603,0.00281423052749119,0.00692742123241419,0.00595109942636762,0.00260922244220696,0,-0.00660726815012469,-0.00341429533432092
"998",0.00107106241494348,-0.00713554203037303,-0.00279093780369288,0.00151133400100978,0.0182372527265016,0.00860472366636045,0.00780816541123852,-0.0097161345488127,0.00291457294543851,0.00761322130876096
"999",0.00241355916627572,0.00268691930355369,0.000932825674877957,-0.00452631575615015,-0.00107309377806186,-0.000106394012836963,0.0114371117989092,0.00510733627940474,0.00678095395188438,0.00906686105773313
"1000",0.00634037082144445,0.00541073021610949,0.0059117804158122,0.014597219347591,0.00697938516049956,0.00213327397874652,0.0109428561950613,0.00909319344211323,0.00155433349452783,0.00636464767940859
"1001",0.00311041839126291,0.00358805484638447,0.00373119464799343,0.00344073570503589,-0.00714394788876238,-0.00276765279406144,0.00696610413528731,0.00715622674858563,-0.00199529992634417,0.00520837720647793
"1002",-0.00143121935464396,0,-0.000929277334719147,-0.00107153487707412,-0.00204018988603694,-0.00352192186352052,-0.00307876489731407,0.00131574727775896,-0.00288781185736087,0.00370098782268258
"1003",0.000398156706499009,-0.00689484572483401,0.00279045201390704,-0.0032182874105976,0.00893115201795958,0.00385579683075266,0.00799255562040435,0.00630755607237488,0.0026733995938395,-0.0018437084596814
"1004",0.00143249050650063,-0.00128583277187244,0.00742109860909435,0.00086112725688392,-0.0195846791354755,-0.0105047010398686,0.00396505782844292,-0.000522279545113413,0.0162938596861544,0.0107130102608699
"1005",0.000715320663352115,0.00926878107851081,0.00920840604244177,0.0128025176148043,0.0169200835254744,0.0112434841928535,0.00448748258332388,0.00966796981499884,0.00357095173028021,0.00036549207135006
"1006",-0.00158836057014966,-0.00459176296734809,-0.00821195970789912,0.0050989197445217,-0.000751405215444589,-0.00203155444974179,0.001250622362309,0.000776653032329433,-0.00493797084768133,-0.0120569444895691
"1007",0.000238648842230127,0.00666336239226251,0.00368002706406712,0.00697498554383214,0.0110639126831964,0.00503500310196281,-0.00124906025961646,0.00672369593558741,0.0123330804373718,0.0188608017722003
"1008",0.0103380679700864,0.00814684838775515,0.0091659903300112,0.00965589853641835,-0.00754359223938139,-0.00309112460374106,0.015546805189284,0.00899024576134511,-0.00519031859003516,0.00435584443840731
"1009",-0.000550923694998651,-0.00202031962901017,0.000908281692594048,0.00457374518988152,0.00117796203451026,0.00235221169458022,-0.0177720518086333,-0.00509140508967754,-0.0235507246376812,-0.0133719597444494
"1010",0.00519780825586791,-0.00632607670756646,-0.00725947582680109,-0.00248318094164723,-0.0220273258807372,-0.0107735115617299,0.00412007030468597,-0.00230323615175432,-0.00282007421150288,0.0106226410499182
"1011",-0.00195889960544027,-0.0114590439517531,0,-0.0105809301581744,0.00437340820179655,0.00517551604975086,-0.00535225435667352,-0.0143625475805887,-0.00401870224077916,-0.013410585848192
"1012",-0.00196252815263143,-0.0054092019670513,0.00365597626670588,-0.00922610591624673,0.00533392592029958,0.00665085487597405,-0.00035891800123844,-0.00312271695235111,-0.00186804151732733,-0.00367371914114689
"1013",-0.0012582767911028,-0.00492151551009479,0,-0.0103708640254304,0.00541367085765221,0.00341071969754236,-0.000358694813580751,-0.0031323325359498,0.00404246887194981,0.0117994381284996
"1014",0.00354396574879301,0.00702757884305316,0.00728602949005097,0.010692864315774,-0.00559908711799229,-0.0039293293631204,-0.00179535024687494,0.00418971943916779,0.00589031486319391,0.0112973335278741
"1015",0.00902452108524399,0.0294651696818202,0.00904178340455131,0.0201018283725107,-0.00779883335179221,-0.00287906145118855,0.00449593169365214,0.0151240286236898,0.00407681405153615,0.0064864718915163
"1016",-0.00163326263122288,0.00477047390941499,-0.000896384918070869,-0.00871203283485567,0.00895073836051519,0.0067361186746755,0.0028643349653712,0.001540957012091,-0.0104090058108441,-0.00143220592840976
"1017",0.0072445503693408,0.00924517375447276,0,0.0029297109414359,-0.00638324320835071,-0.00276100450451389,0.0067830467485388,0.00641177645310775,-0.0101454753417649,0.004661289919627
"1018",0.00170163568546755,0.00990350005443164,0.00269084041909529,-0.00146052575026678,-0.00468120728327714,-0.00244993723002418,0.00939721516065961,0,0.00557684067259268,-0.00107079602915094
"1019",-0.0098057074348521,-0.00833556501093868,-0.00178883779715866,-0.0077310793926656,0.00721993272617083,0.0025618961267988,-0.0119441458563203,-0.00535149465327522,0.00217348433796283,-0.00107179677897651
"1020",-0.00132563769192662,-0.0064277970947878,-0.00896076213419417,-0.01094964900665,-0.0137941426719043,-0.00777328171131952,-0.00213349330359958,-0.0102486053903682,-0.0188453782617007,-0.0100142801895847
"1021",0.00226455314234264,0.0126898027904305,-0.00994546178101163,-0.0104319940950391,0.00792971362992012,0.00332666781899849,0.00391949670409542,-0.000258552713455096,-0.00129571649304228,0.0101155804464559
"1022",0.00568657923685389,0.0100739090784427,0.00639262442895894,0.00774541238028026,0.000436659741051226,0.000107123216876115,0.00496853811312836,0.00699064811799177,-0.00511331759988787,-0.00858361088916537
"1023",0.000542101283670826,-0.00267586023247635,0.00907449584251441,-0.00597794857861222,0.0095019300839323,0.00502747626412914,0.0105950744925807,0.00539994411308542,-0.00199443846276126,-0.0126262752838782
"1024",0.00387110727606244,0.0053657275153578,-0.00179880188006187,0.00880564976571074,-0.0151463195994964,-0.00606606528467446,0.00279603748782953,0.00332485680219419,0.00814756303700692,0.0222871715082313
"1025",0.00246774801171901,0.00558011463477004,0.000900839126991348,-0.00340625887598467,0.00450420144351882,0.00374686106075584,0.0139397909706553,-0.00254919107575624,-0.0246264402370709,-0.00857762194444589
"1026",-0.0174629275298777,-0.0243669366092848,-0.0171014766781417,-0.0316172581419635,0.00524910860310634,0.00458743212242929,-0.0156383348793505,-0.0171222413516489,0.0183694129602125,0.0126171730460689
"1027",0.00751634149985025,0.014095160084499,0.000915581915736707,0.0105890713208565,-0.00761505738472501,-0.00392832627902362,0.0118712578216258,0.00832019875699008,-0.00314709858111084,0.0156639803234693
"1028",0.0160089188650205,0.0246281806476947,0.0201278729754708,0.0242304221349945,-0.00495033304544701,-0.00465028276174961,0.00465841558016011,0.0180509513963176,0.00716106903677027,0.00736068056253858
"1029",-0.00191230535608955,-0.0033317614925642,0.00986567919949755,-0.00745959369500482,0.000221114084126617,-0.00236149573137745,0.000171791842101587,-0.00303950423451016,-0.00267588678877939,0.00974249329415966
"1030",0.00222251774888038,-0.00501469328836901,0.00799288705249346,-0.00128831202737967,-0.00829070205837801,-0.0057051452436705,0.00257544843432655,0.00152404148426588,0.0134151018799946,-0.00654715488960811
"1031",0.00282884102187486,-0.00287941927856117,0,-0.000215039152968499,-0.0101426626646227,-0.00617020783397559,-0.00907721047189103,-0.00608802074750403,-0.00408466726364609,-0.0055498412586894
"1032",0.0062524192498028,0.00601672062435687,-0.000881175411374779,0.00129051242851119,0.0051806358531461,-0.000435207149657613,0.0112342715511495,0.00280732614219614,0.000151822872495266,-0.00279037104622348
"1033",0.00454691446635569,0.00717680187881919,0.00617315736797641,0.000429668528459271,-0.00918616671870764,-0.00686492131909144,0.00256366000387653,0.000763642151814237,0.0110875309660747,0.00664576963206298
"1034",-0.00226327523587677,0.00190044244500465,-0.00701164722392533,-0.022971425658562,0.00870517453328779,0.00570564865518319,0.00238666745952276,-0.00940987814181671,-0.000525702272237361,0.00486435090443704
"1035",0.000378223676722467,-0.0101943674070495,-0.000882322098005983,-0.00944818158633942,-0.0115442614570641,-0.00327311445613809,0.00323128379411597,-0.00744587395496188,-0.00165327262664072,-0.00587820501003333
"1036",0.00597031431174599,-0.00047899922895267,0.000883101277778131,0.0122003568346942,0.0144010056660153,0.00459721384923917,0.00627250648885114,0.000259135046031034,-0.00398945409155649,-0.00347824910264893
"1037",0.00240355939528314,0.000239582964746132,0.0088264150218289,-0.00504051247923776,0.0006698102660192,0.000326319184396295,-0.000168592344113261,0.00206883585615247,0.00476110917980832,0.00488653099623337
"1038",-0.00314758661983605,-0.00167727597839318,-0.00699935282454933,0.0019823224156581,0.00446898526826112,0.00228783795108467,-0.00336993607570235,-0.00567773766932189,0.00767208742396597,-0.0128516878535987
"1039",0.00631552771685273,0.0112794484953975,0.0140968935340076,0.00835343075898143,-0.00322537247653587,-0.00141239012389083,0.0028740187618792,0.0124577495199503,0.000970403814507748,0.00738913410732644
"1040",0.00298845231048284,0.00427140612878651,0.00868818093788182,0.00348804907457079,0.00156205961663325,0.00369943605726419,0.00134877443934611,0.00845954076043709,0.00700959700180781,0.00314354882990564
"1041",0.00208586478092387,0.00472609634698329,-0.000861342143217869,0.00608311907359504,-0.003118933096802,-0.000216606098339178,0.00387201677040316,0.00279607093967082,0.00274001050933093,-0.0010444823480118
"1042",-0.0200702351514984,-0.0275166875115673,-0.0275862859001982,-0.0319585174044522,0.0149734557130463,0.00965172200277786,-0.00905583252993136,-0.0240812335567725,0.00649870005173336,-0.0013942307795789
"1043",-0.0061441236628168,-0.000967233954767166,0.0017731847993343,0.000892147015820077,0.00363366317923242,-0.00247043545207903,-0.00795428435252632,0.00545472750774145,0.0089515156112745,0.0223385505785685
"1044",-0.00068698512571741,0.00145211275358403,-0.00265501803019341,0.0024515894412025,0.00636236605402885,0.00258479455259941,-0.00545868660073412,0.000258471048073972,-0.00749035733729753,-0.00887669868527741
"1045",0.0106926015500082,0.00991066467220936,0.0133098387489559,0.0120054266285816,0.0058862440773999,0.00322095704828729,0.017838843250654,0.0178201023373017,0.00659443893887568,0.0220461048357377
"1046",0.00619681071781186,0.0117282483167185,0.00963214573999904,0.00593134308241949,0.0013001531793333,-0.000427649967481125,0.0208966058103885,0.0134483690518352,0.00203813502554451,0.00168514618857385
"1047",-0.016672970865515,-0.0160870831376146,-0.00173466215041007,-0.0102642738282822,0.00289890402762683,0.00113822538850528,-0.0269066365756959,-0.0160242564643615,0.0172162932669973,0.0151413553204189
"1048",0.00213861911810787,0.00673213432473152,-0.00868787910510804,0.0136803624396857,-0.0153729993997175,-0.0052547831525247,-0.00797300877744878,0.00508942353171626,-0.00078555310137518,0.00397754323492205
"1049",0.0172242082161997,0.0128973253635372,0.00964056138747993,0.0198086385202902,-0.00978571603423817,-0.00679094601049834,0.0143639380006091,0.00860749537193284,-0.0130789167106762,-0.000330205386527171
"1050",-0.00749236177991996,-0.00848870401169954,-0.00694457079699617,0.00106718539264761,0.00832771804412147,0.00716344931172141,-0.00859737097304913,0.000502199843230411,0.00912455671300028,0.00495373116318754
"1051",-0.00785068869844352,-0.00808557879988625,-0.0192305901376388,-0.0140723890068108,-0.00638683261155948,-0.00247828203313594,-0.00646153981067543,-0.00777703320416445,0.00265514879131024,-0.00460062643848858
"1052",0.00875000291650974,-0.000239509233068369,0.00445612498958536,0.0134081999990496,-0.00609518136739573,-0.00237718418011068,0.0124934422434004,0.0022753413565848,-0.00257658171645725,-0.00858377702770841
"1053",-0.00143336330194577,0.000719297335844971,0,0.00192056013271746,0.00970122908431592,0.00584742198858423,0.000507321264602068,0.00327940198714738,0.000358804532442303,0.00399601803386762
"1054",-0.0185057130778572,-0.0230050868642229,-0.0248444569118673,-0.0296059991905143,0.0167860227109249,0.0085052704562063,-0.0155431838080082,-0.0226301980599952,-0.0117638616522814,-0.0162520558719252
"1055",0.0069261937891365,0.00392445841325606,-0.0163784531123174,0.010316091895834,-0.00564774315529437,-0.00234872341340009,0.0113266062075297,0.00102893176457464,0.00326629155066294,-0.00573161612253437
"1056",-0.00603784869629065,-0.00464217084339535,-0.0703056008385818,0.00586573201748442,-0.000437322062669443,0.00224684172154888,-0.00678783671940775,-0.0187612108371432,0.00463029948900107,0.00271274688097622
"1057",-0.0114570806063135,-0.0252822809014642,-0.00198985581438405,-0.0166307293620629,0.0149710587258145,0.00363000093454802,-0.00802983942260604,-0.027501016151701,-0.01865185785214,-0.0365235273160286
"1058",-0.0185127740722061,-0.0307226474717129,-0.0368892224178861,-0.0204259516759282,0.011305433807671,0.0085091815490479,-0.0130900862502404,-0.0250472172730767,-0.000220143825636065,0.00596703307699742
"1059",0.0132350140930948,0.0350741229331366,0.0455485469612613,0.0123318546760607,-0.00766594268157017,-0.00305837147891608,0.00837715425002616,0.0256906977618139,0.00535816187029647,0.0310536687711132
"1060",0.0036371534173627,0.0107930990023966,0.0267329003384578,0.0017719706167878,0.00268276644096166,-0.000634569344890257,0.00882634345165778,0.0237393815031677,0.0102211724449064,0.00575298742614816
"1061",0.0154978527160956,0.0245840816440703,0.0289292297707175,0.019234893627871,-0.00588506051916216,-0.00518792651772204,0.0109797073523792,0.0237968018871118,0.00556481916473284,0.00471070698178733
"1062",-0.0034686473101011,-0.0026658463312822,-0.00374867998493578,0.00303698041679157,0.0033359685225236,0.000532804731973036,-0.00899384144133564,-0.00723142157730972,-0.000646801787025919,0.00736764965761338
"1063",0.00286186994678617,0.000728847527653009,-0.00564453225003458,0.0131919840155588,-0.00128698552178241,-0.00127693078177382,-0.00753417466602235,0.0088448352282684,0.00927718786169329,0.00199472211951734
"1064",0.0095631991174101,0.0150558483343455,0.00189229171322336,0.01152610490883,-0.00751828220489303,-0.00511166760459492,0.00465841558016011,0.0105726039720995,-0.00798058309763683,0.0033178730098975
"1065",0.00305614201184046,-0.00885176440470914,-0.0245515532480585,-0.00105522998698504,-0.00248948096908741,-0.0026757888492992,0.00507558492077731,-0.0109722566769987,0.000287271941622924,0.00264546644963271
"1066",-0.00243724454775185,0.000724175120414339,-0.00193603158814337,-0.00506953130144527,0.0014106427267051,0.000321092335866524,0,-0.00438590662440852,-0.00517019981222888,-0.0135224126400227
"1067",0.00671864988973625,0.00410022549927613,-0.00194001171959379,0.0114647458138388,-0.00769270058700433,-0.00289665572795206,0.00448114764581464,0.00103614723755729,-0.00238188260916128,0.00568367458562014
"1068",0.00690098705583386,0.0100889257470753,0.0155491923207081,0.0128043904902611,0.00797042897812816,0.00344373520280095,0.0116679776052984,0.0111315667067478,0.00332820328993977,-0.00132973490910149
"1069",-0.00135556553516447,-0.00546965991588777,-0.0124402512496353,0.00870481199162931,-0.00205837910353746,-0.00257369370997496,0.00746250385888581,-0.000768368349359227,0.00858154624044927,0.01564586580112
"1070",0.00422360730728255,0.0119561291263703,-0.00193790762195223,0.0160263110170549,0.00486167669190096,0.00213465689425929,0.00235685358572768,0.00922434287003537,-0.00471903328529233,0.006882928416728
"1071",0.000825751138746611,0.0054346079715164,-0.0135925079180407,0.00849347333149941,0.00108477739592505,0.00225867850001427,-0.000839664241641502,-0.00025425862065076,0.00459769406460553,0.00911459275608784
"1072",-0.000149609131376738,0.00258527206394166,-0.0196849178741966,-0.00200504573113747,-0.00400904629745424,-0.00504409661453897,0.00168109005014827,0.000507801373796468,0.0158038262529698,0.00096772869811601
"1073",0.00315209050161025,0.0114863764256454,-0.00903610658100951,0.00542484862919634,-0.0150129774825725,-0.0043153719109521,-0.00134297869419631,0.00736048905693765,0.00232313969046527,0.00290047881931033
"1074",-0.00254383631242883,-0.00370793791497726,-0.0081054299279214,-0.000999347410009066,-0.0019883430471801,0.000108277231436027,-0.0104180543032293,-0.0136053465548969,0.000912979318971052,0.00192792795831886
"1075",-0.00345024932438043,0.00790868919902898,0.0194076188436016,0.00100034710429697,-0.00531255872544156,-0.00292487472244762,-0.00747165801405181,0.0107279333940482,0.00806967258682434,0.0237332348437118
"1076",-0.0030106427788269,-0.00138481025039816,-0.00701415624133539,-0.0117906740885143,0.000890061218655314,0.00130399528647973,-0.00102634435981841,-0.00732878588014707,-0.0071001320590246,-0.0184837784171399
"1077",-0.00747390339890608,-0.00970647782941825,0.00201831746969927,-0.0188070380335835,0.0107831491121637,0.00564247619053049,-0.00205513076486874,-0.00789227008562277,-0.00722096191265387,-0.020427623687187
"1078",-0.0000760679553102328,0.000933344517880297,0.00402815428060643,0.00824426054646432,0.00626884952120332,0.00388439117422279,-0.00120132688861652,0.00307943328113502,0.00204782852872087,0.00782006312591998
"1079",0.00076057411406083,0.00349728272958294,0.00702122066997179,0.00306628405921128,-0.000765286767728912,-0.00333237081655091,0.0135742174421891,0.00818615243658849,0.0134602119856329,0.00258645032519977
"1080",0.00364863754438671,-0.00232327437266466,-0.000996034001490065,0.00122267522249064,0.0135624005747228,0.00733329019925844,0.01101832097238,0.00304477070514664,0.00862252289301879,0.00515972166490997
"1081",-0.0112086539348659,-0.0251512101191927,-0.00299099463048014,-0.0250357405294391,0.00226607918943444,0.00246245588778904,-0.00989281761747174,-0.0146723278218116,0.00606680442467833,-0.00609568631687829
"1082",0.00574431255140628,0.00860001718612513,0.00299996751721565,0.0144049494200398,0.00430658681651774,0.00128162475068461,0.0077898651358026,0.00770257703126376,0,0.000322850943261122
"1083",0.0136317211684158,0.0272383005129797,0.0149552040659724,0.0236677305042854,-0.00643255405076981,-0.00394663307597554,0.0115950502621516,0.0168149223441005,0.0039060304758598,0.0158115350310737
"1084",0.00510909686184013,0.00691745350944095,0.00392945790930943,0.00884585807315075,-0.000862855575438748,0.000749694739493822,0.00714294945705407,0.0107743927765696,0.00163825938566542,0.00730619171549063
"1085",-0.00104659845117083,0.00160293787462651,-0.000978576081577809,-0.00817040775376632,0.00377977278362995,0.00353086712215878,0.00494759529755706,0,0.000885852498096806,-0.00283811777633758
"1086",0.00860506752047518,0.00983032902706782,0.000979534630738632,0.00863947437388535,0.00968238923986342,0.0042647504965645,0.00935536358354172,0.00793260891174485,-0.00333621581453702,-0.000316316289468599
"1087",0.00652893533486143,0.0178856627576578,0.00195667059437943,-0.0017927054119149,-0.0102288774223419,-0.00286658371841031,0.00455288647824936,0.0108213435204141,0.0192648715922641,0.0060107715714699
"1088",0.00324305945768999,0.00400361008587491,0.0263669882965585,-0.0081818209126433,0.00764364301619258,0.00383340015318812,0.0111687581781597,0.00389290401214493,0.00415556308623799,-0.00723270247891861
"1089",0.0023509133965558,0.00443038108906135,0.00190287435120684,0.00603607724150623,0.00309814085079663,0.00201503590842322,-0.00480264630265936,0.00484732732059046,0.0170203436180589,0.0104529163490235
"1090",-0.00153909852795509,-0.00220541969482124,0.00284916538259927,0.000199956541742541,0.00160437514391343,-0.000307734557273509,-0.00016060973327614,0.00144697679294059,-0.0128633659140043,-0.010031372377705
"1091",-0.00359709546853437,-0.00773652289907767,0,-0.0221955693769957,0.00566010998024202,0.00265387804076012,-0.00675663850869779,-0.0093928092534703,-0.00352369513932049,-0.0104496070956075
"1092",-0.00663081514622044,-0.00757418407291444,-0.00189375470261888,-0.0165642693427077,0.00445918294061198,0.00254112209115798,-0.00550726735341878,-0.0111842290332314,-0.0143448687501713,-0.0160000118565692
"1093",-0.00904836094363337,-0.0255891275496397,-0.007590297684687,-0.00956546441779804,0.00951553032419672,0.00496349663771523,-0.00146601348599373,-0.011802152700556,-0.0288363576480433,-0.0669918253132131
"1094",0.00441583165476667,-0.00483740588071691,0.00573646387162552,0.0130167003533308,-0.00439856210378042,0.000525588579489256,-0.00538180934166255,0.00870850735888107,0.0127552937007369,-0.00313697441194594
"1095",0.00387486299798812,0.00555512045980122,0.00380193679636798,0.00186533302894398,-0.00105159939052069,0.0014703000159193,0.00393543510579542,0.00419337347765447,0.0143152233795893,0.036713179193959
"1096",0.00853627712831262,0.0112804943026223,0.00473485282044739,0.0117915040198919,-0.00716001549146916,-0.00482469370965721,0.0138843220302152,0.00245648590767567,0.00352821944876425,0.00910628911108069
"1097",-0.0105248837539279,-0.0168454453168558,-0.0169648643793158,-0.0220812214174856,0.0057264285553853,0.00358323247501224,-0.0111164870716332,-0.0161723556820712,-0.00919540943321462,-0.0320855705109503
"1098",0.00476042710860258,0.00324177980084173,0.0028760647983519,0.00292715873578753,-0.00632722036708744,-0.00220503762144475,-0.00016283529522243,0.00547920265600799,0.000341224255415495,0.00103589746505772
"1099",-0.00769916913682689,-0.0159244250784273,-0.0210324184661549,-0.0218889581873297,0.00902076976999067,0.00389429719318901,-0.00912506100809485,-0.0118898181783776,-0.00654881660546602,0.00172481566061466
"1100",-0.00634137938306267,-0.000468939868672247,-0.0058592836121425,-0.00149175833209736,0.00557418792665443,0.00241061724972624,0.00230218225127032,-0.00200547454739153,-0.00178541503174445,-0.0130854680616797
"1101",-0.00015002799301711,0.00187716257226622,0.000982250721778932,0.00320158208867682,0.0102500888132937,0.00292836573705824,-0.00147640400048277,0.0072843644429248,-0.00433370036230651,0.00244246696417449
"1102",0.00893573414976911,0.00702544099644564,0.00785077780314869,0.0161702146563503,-0.0132517534794044,-0.00573501408498944,0.0111729995633409,0.00798000837924806,0.00594169524866328,0.02018793134022
"1103",0.00238153349299997,0.00837232414580158,-0.0146056315968759,-0.00649087764494194,-0.00041976629912166,0.00104870809159729,0.00194986889310833,0.00569057957810326,0.000343324161676151,-0.00784711418311368
"1104",-0.00794445690193979,-0.0161440442566538,-0.0108695913372827,-0.0080083036605606,0.000524503285509015,0.00240977602264447,-0.0102172449731013,-0.00787223049870933,0.0126331004174296,0.00928471077985238
"1105",-0.0116010805514584,-0.0241444914315502,-0.0149850855705557,-0.0208199700056262,0.00482591871485294,0.00135897900216508,-0.0104865065858575,-0.0176052796936098,0.00230522061478,-0.0160136901516122
"1106",-0.000833045503237706,0.0031229427331243,0.0121704024885467,0.00998043824937489,0.00375863304691992,0.00104330008335962,0.0029803501002057,0.0055534620329678,0.00514099972751136,0.0135042207483271
"1107",0.00333456247448471,0.00933903292775318,0.00200416067562226,0.00214823051318169,-0.0046803528557724,0.000104122015915475,0.00412754777965674,0.00301202662384559,-0.0000672589021404324,0.0181072403749749
"1108",0.00460793773126955,0.00972713817478632,0.00899975779770656,0.0128620132868975,0.00856923838876966,0.00552539794114937,0.0129892875258399,0.00725721866601825,-0.00242294383600838,0.00369129388523048
"1109",0.00383443374410741,0.00798887292519312,0,0.0105818673084028,-0.000414455226153132,-0.000103255310902606,0.00178540337242206,0.0111800448327988,0.00998513014448021,0.00568367458562014
"1110",0.0104111819965975,0.0219113620156455,0.0178396004296768,0.0163348840889042,0.00228029807617092,0.00155556634815968,0.0174984273821994,0.0122850947618356,-0.000400788251184836,0.00565158721344039
"1111",-0.0224610258433859,-0.0278284684496696,-0.0126581764643997,-0.0179271148431203,0.0135146635102645,0.00824024180594574,-0.0281848305188405,-0.0177185002537831,0.00180436381852678,-0.0125619145801649
"1112",-0.00106174832622208,0.00821223626064316,0.000985982793067164,0.00944199528395639,-0.0190493401014494,-0.00597053395953584,-0.00573469731130183,0.007165881858469,-0.00273500092762313,0.00870430105841091
"1113",-0.00994440324721169,0.00744684886581859,-0.00886695828912032,-0.00498859457119549,0.0057424289139838,0.00393561323955738,0.00362555656422558,0.00147159317722045,0.00481606020066883,0.00398275562528294
"1114",-0.0105814526919037,-0.0157080400245176,-0.00994033862932375,-0.0160851863565665,-0.00757831476144821,-0.000618712341947325,-0.0142859013545747,-0.0100440805935313,0.00173076153820562,-0.0115702605873167
"1115",-0.000619559880307152,0.00938746258080858,0.00803230466745508,0.00785551789345917,0.00460283059643873,0.00185782524129441,0.0119942373522484,0.00296969895929933,-0.00039871080273024,0.00936459327804839
"1116",-0.00418753508641312,-0.0169729318630751,-0.000996034001490065,-0.00716244882786965,0.00780908108826917,0.00216350055174397,-0.0047739840510127,-0.00764894188750831,-0.00405531184756425,0.00828362085452339
"1117",0.00763107828240783,0.0130087226140259,0.00697907406370968,0.0078508019740835,-0.00402967775457808,-0.0040092067577987,-0.00926240699872483,0.00372977862616342,0.00500634143256584,0.00558665132076031
"1118",-0.0139102820070212,-0.0263832291115101,-0.00990096909755545,-0.0216841763456169,0.00767646665318633,0.00319995003129603,-0.0237058029280189,-0.0173392805522432,-0.00876722248628092,-0.010457541356911
"1119",0.000783862589043283,0.00263774852166376,0,-0.00172166303867116,-0.00504387342779444,-0.00216077710741136,0.00188086755485162,0.00252084506541439,-0.00984991256198364,-0.00660506552415063
"1120",0.0126858688449412,0.0141114533035773,0.019999986103622,0.0150894529840728,-0.0151060539767836,-0.00794032420143809,0.0157019507606189,0.014583778355199,0.0060905053504634,0.00698149320234909
"1121",-0.0177855904171516,-0.0360847820494319,-0.0196078297804899,-0.0214480667383177,0.0181742256931599,0.0108099741374295,-0.0164673676206976,-0.0195785727130225,0.00302681782507319,-0.0267415394978376
"1122",0.00220465365076494,-0.000489601589313549,-0.00300017017273246,-0.00759578437576225,0.00453984160450549,0.00277638005328074,0.00700475084839125,0.000505170212192985,-0.00100586108522871,-0.00407053551353975
"1123",0.00298402397540176,0.0124848407259399,0.00300919827965496,0.00131216233341558,-0.00472488201971766,-0.000717639372510015,0.00848310870592694,0.00319174926448129,0.00651138479887625,-0.00442780233597684
"1124",0.00511602903392538,-0.00362674958240083,0.000999902320041102,-0.00152859810613448,0.00123818502035977,-0.00153881951023294,0.0105991258961307,-0.00254516376373692,0.000600220080029246,-0.00547389412708488
"1125",0.0137042255564421,0.023268356752534,0.0169831528955764,0.0183726136539146,-0.00443197945396023,-0.00133669686520166,0.00882298861314834,0.0130136486618602,0.00486566689905787,0.000688055927610343
"1126",-0.00602553361054792,-0.0126058245569975,-0.00118920050325444,-0.00995686419982011,0.000621379670626032,-0.000411746946021863,-0.00214513730247434,-0.00881631126418436,0.00152566998957515,0.00446882846379237
"1127",-0.00287561279149295,-0.0122758822777612,-0.00198418031403391,-0.00131447792026018,0.0076565020443824,0.00525072314530961,-0.018356185533613,-0.00304956362922582,-0.0175508902062754,-0.021218265704642
"1128",-0.0116132045434741,-0.015660184952209,0.00596426122081617,-0.00175527806941889,-0.00421004742918796,0.00419972947511638,-0.00108810454341801,-0.00994128878434286,-0.0140218488343495,-0.0118882007975992
"1129",0.00891082590125003,0.0111112010930867,-0.00494051815345331,0.0116482996304228,-0.0137136655132986,-0.00387608165156172,0.00527615523295855,0.0043768921897096,-0.00362367713741552,-0.000353779382827213
"1130",0.0130527597275349,0.0119877730667293,0.0119162179561645,0.0136868139232353,-0.00805044093422769,-0.00921474642348163,0.008295099850677,0.0125608655316196,0.00349968444382576,0.0176990911858448
"1131",0.00856414559121688,0.0194968171969947,0.0157019522503108,0.00921544021879805,-0.00664041991891351,-0.00599335935337175,0.0110810701978643,0.00911426647352842,0.00642770765769596,0.0180869597716493
"1132",0.00956244028263975,0.0186395402749577,0.0077293705126138,0.0108304122607257,-0.00159195765881859,-0.00343143650490629,0.00132808616222468,0.0130455728260892,-0.00801734648811947,-0.0105910798016576
"1133",0.0147762259104471,0.00879270252605791,0.00862906297534383,0.0117647447970159,-0.00159901028269305,-0.0024990309214229,0.0179107488741082,0.00841985589597716,-0.00732881506849314,0.0013812676985363
"1134",-0.000821685405087758,-0.00777390673119005,0.00190108243814024,-0.000415273945415739,0.00224266928642591,0.00629053265599677,0.00619083789816255,-0.00736742558606673,0.0186297669937789,0.0134482335920072
"1135",0.00119601569936356,-0.0104461849659895,0.00569253446459528,-0.00664721841236771,0.00511524659548823,0.00177068580188289,0.00615292557724101,-0.00395852453992651,0.00867031739245672,-0.000340247139329009
"1136",0.010375213021858,0.00791709086266801,0.00660382929499281,0.0138017262500372,-0.00296854168906135,-0.0038475805687348,0.0125521716556201,0.00596119032460019,0.00161164457426244,0.0211027479228436
"1137",-0.00709200942236787,-0.0147579933494356,-0.00843496937906552,-0.0113450251687184,0.0141429198050596,0.0106487090955034,-0.00349635675276316,-0.00691325114022989,0.00737516623701651,-0.000999986380040063
"1138",-0.0180804333007594,-0.0374487355632307,-0.0122871366012334,-0.0279573486178677,0.0149951591955586,0.00764366118606197,-0.0188197965575053,-0.023620196735344,0.00891844259567387,-0.00767430506191968
"1139",-0.00431911857958855,-0.00803207575528686,0.00287046445194217,-0.0100881062132717,0.00340832706650884,0.00143508151287275,0.0034137160540999,-0.00127326981255071,0.0077842076069452,0.00874238413852768
"1140",0.0033485289226971,0.0156879929317106,0.0190841577183118,0.0162620135150546,0.00277974918676738,0.00163740000718793,-0.00842404925730544,0.0104539874238967,0.00896769630247563,0.0136667549848453
"1141",-0.00690239049249108,-0.00722474745085999,-0.00936333276783263,-0.0106677930545386,-0.0142710177171772,-0.00572328628541241,-0.0111092114700363,-0.00782254441565911,0.00259500455816153,-0.00559029126745914
"1142",0.00580479813978441,0.00150576541052416,0.00756153184877251,0.00625409791194675,0.00166637351357291,0.00411209768647947,0.0109035889856406,0.0050865633551096,0.0042707650439715,0.00892861944212275
"1143",-0.0082010154914508,-0.0175393829032303,-0.012195220452093,-0.0115732324459762,-0.00967021095944109,-0.000614882575282527,-0.00898824421582101,-0.0129049808771226,0.00882738419125095,-0.00557203579296839
"1144",0.0162312475064681,0.013261803705414,0.0123457799603628,0.0145275735175312,0.0207894915150819,0.00379075322605948,0.01731545885135,0.0115354042449038,-0.0121990350297424,0.00692156308141456
"1145",-0.000602699341968993,0.0135917863134498,0.0103189974824847,0.00299187694902336,-0.0118286340996969,-0.00489841228456656,0.00745659031824308,0.0060823639742944,0.00879348225026555,0.00327327776015629
"1146",0.0138713392586749,0.0273154752217561,0.00835654336295133,0.0159812322476318,-0.00770297195368064,-0.00553736234274493,0.00643601347967238,0.0118384754342795,-0.00762723990187819,-0.00489389755420977
"1147",0.000669272667577658,0.000483780140561718,0.00184166997740198,-0.000629081064465908,0.00755295453080951,0.0038152185816378,0.00511564716169999,-0.000995536580708389,0.00833167334067442,0.00819671052420667
"1148",-0.00557281007110488,-0.00579858747604145,-0.00367664806566648,-0.00209864361516776,-0.0109315918064644,-0.00318434459694095,-0.011293042777001,-0.00647890184018785,0.00781450832098751,-0.00487801563658707
"1149",-0.00373630474524789,0.00680408020364176,0.00184514755977849,0.00336503809614208,0.00684211684404845,0.00422518944317618,0,0.00476543132273055,0.00273298595990812,0.00784313079179988
"1150",-0.0204756278213486,-0.0263091952403322,-0.0165746862359859,-0.0176065650105628,0.000104109347096593,-0.00164245342954339,-0.0268661065561389,-0.0154768061467655,-0.00367625014448247,-0.00680941221417808
"1151",-0.00290952369550002,-0.00421442229673985,-0.00187260205799467,0.000853483962409918,0.00376344936786799,0.00195334985466888,-0.00148801415376243,0,0.000827056418003069,-0.00326472866915961
"1152",-0.00683466393422516,-0.00199110833499383,0.00469032857365881,0.00426342204434738,0.0197873614088344,0.0121053018310073,0.000497032609328318,0.000253699489296544,0.00616568749580604,-0.00818865621833109
"1153",-0.00425269638029857,-0.016463039969866,-0.00933707856948529,-0.00084885528527745,0.0100924760584507,0.00363744464514859,-0.0132385811171862,-0.00481624511618195,-0.00360093515197779,0
"1154",-0.0255471985163724,-0.0304338363178178,-0.00848237299129073,-0.0308052918460577,0.0300269807148446,0.00921220401420175,-0.0293479296852704,-0.0191034316413304,0.0240933488201032,0
"1155",0.00541852829028411,0.00706272238779238,0.00190108243814024,-0.00350729378792081,0.00196945895323419,0.00080231868797398,-0.00621948070653189,0.0111656845670896,-0.000185729316846794,-0.014861261469488
"1156",-0.0468415489315102,-0.0727272212342204,-0.0607211391418988,-0.0571930829228079,0.0355807438775375,0.0132303924069503,-0.0483309396800817,-0.06060582749689,-0.0052635207980829,-0.0378813261809202
"1157",-0.00149649726657475,0.0240895817848013,0.00909090724606343,-0.00653287660814927,-0.0288530155720829,-0.0115737029595531,-0.020643073016651,-0.0032804466319043,0.00690986682588313,0.00418112739105347
"1158",-0.065123570452394,-0.0820570123974501,-0.0480479330447384,-0.0833728603073269,0.0315668592616944,0.0159124148703542,-0.085058787572338,-0.0811851074269598,0.0331993508500772,-0.0371269529125423
"1159",0.0464995580051517,0.0694277232257374,0.0515247177170461,0.0586729655249294,0.00303205349107616,0.00581258128224005,0.0925585542769012,0.0800001760268474,0.00891578533137238,0.00972978201500774
"1160",-0.0441777684856008,-0.0696571991621485,-0.0460001698497129,-0.0530009759174319,0.0297536390150952,0.0132216955335045,-0.0235118348531859,-0.0527915301138158,0.0354071583215281,0.00428252295001075
"1161",0.0448834346610443,0.048817021620561,0.0377359035491276,0.0552010061426156,-0.0504499983088923,-0.0146926296443122,0.0466273921613214,0.0469797453732042,-0.0219383775697288,0.0216773984576242
"1162",0.00673332446107411,0.0251286647503308,-0.00909093623649715,-0.000484689039714103,0.0198036128741577,0.00696571835985593,-0.001460843149376,0.00780389864045361,-0.00456807613469989,-0.00139135691917081
"1163",0.0211650113390052,0.0239551653465975,0.0122326283018299,0.0232614448168864,-0.0101352107420943,-0.0037021194143948,0.0356555953874809,0.0210174059236585,0.0107666175750627,0.0121908874330814
"1164",-0.008539233924999,-0.0174100824313808,-0.00805661003568603,-0.00852474394546665,0.0165548930641866,0.00459587228849268,-0.003707567714333,-0.00839639764550837,0.0123399008322485,0
"1165",0.000668920968205811,0.00664447485273034,0.00101538689349612,0.00716497595169008,0.0175088555831013,0.00700815422892931,0.00124044684290525,0.00655586070025493,0.00287488503765965,0.00860291493408494
"1166",-0.0431185592082095,-0.0539054639712606,-0.0344828670230404,-0.0471894790841524,0.020538312642552,0.00522017009203535,-0.0430091268549873,-0.0331074635016801,0.0189198660580194,-0.0245650104809031
"1167",-0.0163307153220639,-0.0200579922385654,-0.00945365889541538,-0.012444433144035,0.00806865624268682,0.00105792094452539,-0.0199741601606612,-0.0117876972339348,0.0125478054661952,0.0178383776501641
"1168",0.000799267504768553,0.0115690962027457,0.00212082580451778,-0.00100789270096968,-0.00251832278754294,-0.00182462248021098,0.00188712134516056,0.0036919977347718,0.025784935133953,0.00171818966189541
"1169",0.0329104097738679,0.0340177915627853,0.0190477353248888,0.0350656338505093,-0.0137937084007113,-0.00404213575936663,0.0246752648273123,0.0271648931822097,-0.0374884779779724,0.0102917024523768
"1170",0.0140845887248111,0.00425406610530299,-0.0114228086732449,-0.00974914593582077,-0.0284304842011114,-0.0107256824321386,0.0112134213722317,-0.00110201756877049,-0.033883064489031,-0.0101868622966957
"1171",-0.0152441597459863,-0.0276760515469363,-0.0136553319674453,-0.0194437223257118,0.0108205977610896,0.00615324990551835,-0.0210872849092033,-0.017098667997219,0.00413636484018753,0.0044597718600301
"1172",0.0145341101112761,0.0116181493531595,0.021299090926902,0.0170684399258203,0.00986670832790182,0.00320360075711701,0.0148560193695686,0.0134677838143777,0.029647249769974,0.0112705134484055
"1173",0.0287360661016993,0.0267008501465476,0.0135558978137826,0.0323295275883317,-0.0138261862869127,-0.00658000178617968,0.0318391245499756,0.0271317497918344,-0.0201724346640422,0.00337722592734591
"1174",0.00263683612679277,-0.00782967652843281,-0.00411510045154917,0.00143443438424518,0.0160762195795559,0.00691574731593469,0.00390143187193503,0,0.0299615103223965,0.0134635385750419
"1175",0.00443768447802562,0.01944739178771,0.0175617256936811,0.0205300588284778,-0.0154536885109251,-0.00357920767968312,0.0107753917503457,0.0150948893297764,-0.00770522028904908,0.00166055506291896
"1176",-0.0104727605916252,-0.0102295294945577,-0.0091370542993352,-0.00537992280072097,0.0211978747623627,0.00796924281791234,-0.016777438554536,-0.00929404495574737,0.000843990542178652,-0.00696293982860552
"1177",-0.0255499902231768,-0.0270947793953504,-0.0163934136987397,-0.0225777106262481,0.0324861851289406,0.00917100086014466,-0.0241734440104941,-0.0144733066702829,0.0301906457016543,-0.0053421641792456
"1178",-0.0072973567645549,-0.0422051386666875,-0.0218748561236467,-0.0103467664955715,0.0103989949550596,0.00133860753428294,-0.00218557508905326,-0.0190373723470819,-0.00185555004760019,-0.00335688875632811
"1179",0.0282075407395641,0.0305756100419607,0.0191689862182767,0.0296621486805764,-0.0190884447249154,-0.00534923137493482,0.0335886129611409,0.0202383826720653,-0.0318206243352855,0.00909395082323083
"1180",-0.0103916305689398,-0.0206517231285799,-0.0125389249133422,-0.0221961307888237,0.00896765447855197,0.0048977276188864,-0.00724131833535513,-0.0187497855806646,0.0267110681419576,-0.00667547638088173
"1181",-0.0262093452212897,-0.0380158716128733,-0.0232803190551093,-0.0338079832378504,0.0106656270323386,0.00487428485777563,-0.0281086791658683,-0.0288007859426752,-0.00610528030477187,-0.0157930705888282
"1182",0.00646981042314421,-0.0101883223583247,0.00975080886193846,-0.0019995193006842,0.00105521827022459,-0.00304338652775615,0.00311196428175387,-0.00228133644618989,-0.0223021531096097,-0.0023899317720053
"1183",0.00917113621481125,0.00842159401424514,0.0171673481398888,0.00150268919148289,-0.0142316093064826,-0.00295726854892731,0.000912395349075057,-0.00342938104313495,0.0105846777674159,-0.00308004014999508
"1184",0.01384401302803,0.0238169133263189,0.00421928000795857,-0.00275093183946484,0.00846647581479942,0.000573900531291027,0.0056518903712941,-0.00372835588347875,-0.0074492329570105,-0.00480608216168577
"1185",0.0172573799075624,0.0259819762392925,0.0115547969075782,0.0145436678622164,-0.0152882625747884,-0.00745909894518471,0.0193978674935487,0.0146804891672545,-0.0158569656847878,0.00413940847517402
"1186",0.00591847039986826,-0.00294454585329473,0.0103840463948299,0.00172992017473672,0.00726927778574771,0.00192727589661668,0.00818053802439711,0.0000858685274540694,0.00934635926650329,-0.00446586426941942
"1187",-0.00995723907650437,-0.0318962465873753,-0.0143885221009118,-0.029607399260973,0.019066065486776,0.00817371882609441,-0.0197563250573627,-0.0234690121976671,-0.0154519173746062,-0.0169082305750911
"1188",-0.00116345893394976,0.00671152259306584,-0.00104255648161067,-0.00737332514995159,0.00419655243366512,0.00133529471103788,-0.00287910513486955,-0.00175817429410041,0.014251924461969,-0.00175497785306811
"1189",-0.0294584380578583,-0.0300002110760997,-0.0125261911009741,-0.0371418599296489,0.0330839672938981,0.00428627519805502,-0.0478255384816378,-0.025836780528384,-0.0124587723999247,-0.014767839573728
"1190",-0.0323244028129398,-0.0390501088542338,-0.0158562828078351,-0.0702311831279868,0.0375861743358277,0.00929564180933085,-0.0252083696437384,-0.0334536656765928,-0.0261535405531089,-0.0353319713791268
"1191",0.00602510598921446,0.0117033927232093,0.00322241272673307,0.0266096215917793,-0.0185997559315523,-0.00827007861051177,0.0080383484103117,0.00904235910961448,-0.054717538218559,-0.0177581084843996
"1192",0.0237804172698552,0.0285988908707724,0.0053533549517335,0.0150498241804933,-0.0160556705840024,-0.0041690915809196,0.0126730094387375,0.0117430569885866,-0.0138923714538353,0.00338990068006195
"1193",0.0111833858087964,0.0296784177516356,0.0159742417827018,0.0318507792194807,-0.015308103799797,-0.00666098199166165,0.0105890571307519,0.0186317450920022,0.0193552669202277,0.0168919313092548
"1194",-0.0204185885641753,-0.018203920147383,0,-0.0300691488271239,-0.000341665516336964,0.000191659305425196,-0.0249571723731633,-0.0194904725425739,-0.0274544223540304,-0.0269472233298083
"1195",0.00790351992755145,0.0222496256105014,0.0178198107852805,0.013717404931886,0.00692110473704632,0,0.0148496743659616,0.0149846373633908,0.00947379330768272,0.0117601987558278
"1196",-0.0249890464246934,-0.0365779705657897,-0.0257466201507265,-0.0500678088725617,0.0251188076549815,0.00632128740932747,-0.0263767014676235,-0.0343476622110056,0.00228282185699724,-0.0344957184688444
"1197",-0.0284578311402417,-0.0313773487719716,-0.0158562828078351,-0.0210825026107055,0.0275202154192331,0.00925996669559659,-0.0470634543934156,-0.0190325288776177,0.0183475201612997,-0.00504847487959281
"1198",0.021922866386533,0.0223517129764317,0.0128894659411198,0.0154250184219995,-0.0126811520781553,-0.00510239659968859,0.0377671713953514,0.0104961416914857,-0.0206262913495028,-0.001951653922452
"1199",0.0185153176436466,0.0186947333303038,-0.00424177335039622,0.023215793931284,-0.00719824553358439,-0.00417907161617437,-0.007598271051248,0.0062952876835114,0.0115453438946038,0.0140790482234632
"1200",0.0180913519474284,0.0339034900469624,0.00425984263737234,0.0330532528238641,-0.0184576231549061,-0.00696239127619647,0.0276041671669629,0.0272128073448878,0.00645928731208456,0.0208252518572627
"1201",-0.00669584654579924,-0.00842364622700331,-0.00530226234100539,-0.0119308303515084,-0.00738765634689631,-0.00518637623092333,-0.028235309073893,-0.00243601289071427,-0.00816257685330624,-0.00453344997004712
"1202",0.0334455328850487,0.0445992424107975,0.0255864277962827,0.0447310838894011,-0.0141240535478516,-0.0105237658016495,0.0482244103251559,0.0335775642826235,0.0256942529203403,0.0223909381486429
"1203",0.00100340046754921,0.000290647473973227,-0.00831623061510023,0.000525463694717621,-0.00334564947859517,0.00331745664266481,-0.0184793863850748,-0.00797407194026623,-0.00716603155102513,0.00742391804903431
"1204",0.00877226519237384,0.0223577090418623,0.0062893573707401,0.0280914850263596,-0.014546117452233,-0.00340310093862006,0.016277724870067,0.0214351015805532,0.00715600837177011,0.00184234981324116
"1205",-0.00198771750257876,-0.00198807693040537,0,-0.00893793824138611,0.00995745659172709,0.0040005595762922,-0.00694714175614097,0.00466301297797789,-0.00588014228470357,0.00220658761071491
"1206",0.0170939005293802,0.0133750394800765,0.00208350897459586,0.0200979710084426,-0.0145295198630859,-0.00495687726221283,0.0231249827621649,0.0165362849259998,0.00677751681865324,0.0227523610500662
"1207",-0.0190910469975285,-0.0292051276453844,-0.00415799597064914,-0.0338468518147245,0.0172881495500479,0.00654456546269899,-0.0229822661776159,-0.0231163078567563,-0.00477355586683803,-0.0143524120639776
"1208",0.0195459925358832,0.0161989840077379,0.00939444859357086,0.0266667835571976,-0.00621116758167406,-0.00106723565203093,0.0330483215946458,0.00964053804971843,-0.00479645199841494,0.00546057776377684
"1209",-0.0118292530329969,-0.0170794534139643,-0.0155119378762678,-0.01909873897376,-0.000346991538828001,0.00155396593316426,-0.0124200062398646,-0.0144674636226485,-0.0121725225450452,-0.019551117232251
"1210",0.00437578290411889,-0.000868711191681637,-0.0031514507635183,-0.0192107843886713,-0.00712085573440369,-0.00203691633620795,0.00609751824581095,-0.00411066657575765,-0.013135616849178,-0.00147700870732781
"1211",0.0189869779018523,0.0315941239323667,0.0105375722057368,0.0285865461535773,-0.0105819992890364,-0.00184621059248224,0.0295459323780669,0.0250593152901815,0.0110920958080218,0.00517744365051964
"1212",0.0122612819061483,0.0126439003868388,0.0104274502523896,0.0391145959368775,0.00167940192212646,-0.000487251694282542,0.0264894935700564,0.0132295500319464,0.00940320939309913,0.0158204292876116
"1213",-0.019443815841979,-0.0174804823164756,-0.0144476820988056,-0.0198117167938078,0.0254146734854082,0.00857284097632149,-0.0154123306798433,-0.0218563946772422,0.0283815171188295,0.0032597558763543
"1214",0.0101583146887829,0.0180740895736806,0.00209393631205934,0.018444105860016,-0.0174695632347737,-0.00734094022610809,0.00928321616384364,0.00783532289718214,0.0109305999379332,-0.00577620555844283
"1215",0.0348350942898852,0.0590845862379499,0.0386627997818878,0.0607784842139563,-0.0338973590474645,-0.0120657094128516,0.0427411481012132,0.045781391011398,0.0128435428737232,0.0265069102104287
"1216",-0.000233127673750166,-0.012571910428561,0.00402413720052808,-0.00841888523715784,0.0105169312332727,0.00600775710876289,0.00311324679017977,-0.000825945516954807,0.000412810373114469,-0.0042447971617956
"1217",-0.0241057597954931,-0.0498676164839008,-0.058116294706786,-0.0375001994896522,0.0396555610307243,0.0134130803119226,-0.0131036479729688,-0.0338932580859892,-0.0134418056078823,-0.0152752847674487
"1218",-0.0278884384939125,-0.0424342981948428,-0.0127658119303212,-0.0242584179671652,0.0334740385647829,0.0119940208194032,-0.0337174779768603,-0.019966079008732,0.000239088089855066,-0.0119047844473724
"1219",0.0163115761969983,0.0134108408469942,0.00323261304913869,0.0306376339685102,-0.0124734785356734,-0.00239108484773609,0.0202496285168261,0.00407468658806054,0.0100369993417075,0.00620655986768326
"1220",0.0182271214424163,0.0322209605152979,0.00751886027025916,0.0102338861452271,-0.0137333895877632,-0.00469875452608115,0.011341040252584,0.0133331326883015,0.0157340768453103,0.0123368135976034
"1221",-0.00609880405222407,-0.0167224088637601,-0.00213246749535301,-0.0065122850080469,0.00120314941216848,0.00298683298456015,-0.00753453410672122,-0.0051487229521977,-0.00506635799518773,0.00322572541378996
"1222",0.00621613233268126,0.00113410687438353,0.00854720929769748,0.00849721081592114,0.00635293256659053,0.00115222075588095,0.00247202888316678,0.00373810949919862,0.0241731920103063,0.0146481467086375
"1223",0.0128304593368125,0.0181198878908864,-0.00423728040599081,0.0117959673665695,-0.0127964522690361,-0.00450854551794722,0.011975565829017,0.0117441873149811,-0.00828664437733784,0.00492958259453546
"1224",-0.0369094071076762,-0.0631256576893618,-0.0180849663883224,-0.0585300297203237,0.0207397484973204,0.00886649287575669,-0.0449004926151813,-0.0450169557941744,-0.0084134847485362,-0.0220743406300569
"1225",0.00941856547409881,0.0175125571083994,-0.00108356140610921,0.00657108030317,-0.0148998927648719,-0.00487203326344443,0.000911193289677925,0.00326124128922811,-0.00540482339842074,-0.0010748689279797
"1226",0.0188221646979039,0.030630036551083,0.0108461227080201,0.024102335974191,-0.00610184781044287,-0.00460778284035257,0.0258509042203727,0.0260047538683228,0.0164777843664707,0.00968441420898558
"1227",-0.00947400416217681,-0.0209452009080492,-0.00429183703497238,-0.013728782650488,0.0160830395202474,0.00626830484434748,-0.0200533976679816,-0.0207373390518358,-0.00436887772716632,-0.0106571575633633
"1228",0.00494152333871156,-0.00578212799028122,0,0.00621426084491628,-0.00136130275173663,-0.00134125707366106,0.00869261604317439,0,0.000923810639557932,0.00718126704142441
"1229",-0.0158626747987083,-0.0180284912110713,-0.0183191921396191,-0.026926982225618,0.00911797595521335,0.00364628610527196,-0.00951521569573965,-0.0267645449967461,-0.0106714697123242,-0.00249550960909894
"1230",-0.0158769735943447,-0.0106604319183912,0.00109761416045773,-0.0253869753844794,0.0080223982515859,0.00200823395001692,-0.0179442400148448,-0.0163193478687013,-0.0257127230398438,-0.0232309291562415
"1231",-0.0010645661908727,0.00329250223066424,0.0043863667053925,0.00390684325443313,-0.000251294974377259,-0.00372184002856313,0.00719778916643077,0.00614438656585259,0.00311184309592405,-0.00146353550983858
"1232",-0.0190192245146703,-0.0256563490143351,-0.0196512723668243,-0.0321741255405037,0.0059494683765986,0.00277802083946832,-0.0263881193470709,-0.0262594139590391,-0.0245793767026421,-0.00732866692535983
"1233",-0.00392793543008796,-0.00979793299897713,0.007795424597002,0.00348524849771525,0.0111615838143659,0.00305657104803969,-0.00282331163710614,0.00689867185468795,0.0110703241590215,0.00664450312592546
"1234",-0.0220656204035405,-0.0303029533759526,-0.0232043314777461,-0.0323267728544029,0.00980331253853017,0.00342823247273083,-0.0294448860472055,-0.0277172307931967,-0.00290361143189899,-0.0150348950280789
"1235",-0.0018877594546145,-0.00510213013964012,0,-0.0033133837661683,-0.0145212445012344,-0.00635875917154105,0.00350094964623349,-0.000640529606707463,-0.00867565359854827,-0.00819058292561925
"1236",0.0289669509843622,0.0503206608207667,0.0282808315503995,0.0479228342358173,-0.000497051764824286,0.0000952904679158983,0.0244179298696643,0.0326924812016216,0.0197675099057839,0.012387333873749
"1237",0.00284023913986853,0.00640808185321373,0.00440017807583382,-0.00449398142182245,-0.00819894229035378,-0.0019098542772118,-0.00283760422118162,0.00682782071240529,0.0015003300275962,0.0129774726077585
"1238",0.0411497812307329,0.0527594560236997,0.0328587718399855,0.0624004927082,-0.0156159423566443,-0.00583675391035876,0.0461013870289002,0.0554870834485715,0.0194750713244525,0.0117129078004778
"1239",-0.000160067352790283,-0.00576055245972518,-0.0137858090417977,-0.00299945919073985,-0.00501730250535903,-0.000289111982191725,-0.0101559216518907,-0.0175232071339615,-0.00293892896787962,-0.00361785859813823
"1240",-0.00088040273176726,-0.00144829636958244,0.00322590829218994,-0.00300815157916656,0.0140165560272745,0.00443700334734087,0.00164920318916995,-0.00356753746069138,0.00112009664799562,0.00871458986637008
"1241",0.0108921612463084,0.010443982091799,0.00750249522288549,0.0163440378365052,-0.0020230697258754,-0.000576004971602595,0.00932858602039799,0.0137235491982675,-0.0147214691847233,-0.00539956831462385
"1242",0.000317164785908375,-0.000574213811206703,-0.0117024268128887,-0.0136071743053483,-0.0095432754531648,-0.00259455762657934,-0.000725080355214902,-0.00706331596170895,0.00513976789398529,0.00542888193349578
"1243",0.00372239533764285,0.0066071975282127,0.0139936899598043,0.00401299075415307,0.00358127878286818,0.00452806706615427,0.00943066100640588,0.00533484848024135,0.00725413872505043,-0.00863930189363515
"1244",-0.0219365490158754,-0.0342466804055748,-0.0244162016032691,-0.0359729195391156,0.0124904096405347,0.00508255048829676,-0.0238952255261813,-0.0341979140722791,-0.0201888909157812,-0.0127087255023969
"1245",0.0169423138436147,0.0257094522084074,0.0228511536225338,0.0202123264768743,-0.0205605571635171,-0.00686987270788109,0.0198788983597067,0.0149574770541212,0.00253041336378867,0.00367777219365739
"1246",-0.0145974822385259,-0.0342842273410426,-0.0170214591409811,-0.0375919847856779,0.011139022991393,0.003458398851647,-0.017866808396421,-0.031579148142256,-0.0265023386959977,-0.0128252236904338
"1247",-0.00933880687980793,-0.0167064117643142,-0.00432887295767659,-0.00923723625875261,0.0093210732716158,0.00459634936414899,-0.00882039833845483,-0.0102485531062574,-0.021853249526105,0.00408313009436156
"1248",-0.010646087659217,-0.0109225700369922,-0.0108693275156944,-0.0143847151799757,0.0188898510555053,0.00419347810397452,0.00574702571949826,-0.0128647318804186,-0.0350899217751327,-0.0354898435017028
"1249",0.00361421243666427,0.00429476628357617,-0.00219808161287094,0.00648648451990286,-0.00370739718233437,-0.000853503913127329,0.0136405015954115,0.00985397647808917,-0.00366274448075565,-0.00498276289883115
"1250",0.00148271619606577,-0.00763588869252729,-0.00330394320961391,0.00751883776014362,0.0116612214026299,0.00484405940445298,0.00836530360887844,-0.00331903371923381,0.0190375760646284,0.00808941651852191
"1251",-0.0106918079204776,-0.00447568431570322,-0.0143645680310085,-0.0258528322586505,0.0126715601144876,0.00340315148634551,-0.00973851400501391,-0.0150498678436242,-0.00231914584343618,-0.00458549768908145
"1252",0.030260079940627,0.0384012889783405,0.0256408655886358,0.0419024577295903,-0.0249455117031299,-0.00904471100144078,0.0302312287792559,0.0367360777912562,0.0136243369801878,0.0230327116103957
"1253",0.00193656946629628,-0.00541171286194719,-0.00995574353675388,0.0031813047673428,-0.0139100040181229,-0.00323228367538053,0.00141411904844913,-0.0119161410342137,0.00114669387556865,0.00712943567986613
"1254",0.00885892867318816,0.0120918737250855,0.0067039575247978,0.0132137257740863,0.00419882410914729,0.00124039521528596,0.0136809776344868,0.0111078967475051,-0.00712656510240339,0.00111779615846253
"1255",0.00894061765764054,0.00567498426534918,0.00776911021545001,0.00391227725239118,-0.0111206951977629,-0.00409729751413379,0.00492703974030095,0.00784669031194141,0.00173035767823948,0.00483808137586306
"1256",0.000791218034004837,-0.0026729634433541,-0.0121143357725916,-0.00961295067810497,0.00475039515135744,0.000566394041692009,0.00227644814043804,-0.00654019164140374,-0.00895652241003819,0.00444445986150788
"1257",-0.0131234830822295,-0.0157832368340466,-0.0122633668093072,-0.0167891918925264,0.0184887367873572,0.00632091984438676,-0.0108316587290754,-0.0163009189556614,-0.0250468329985969,-0.0117995140293872
"1258",0.0103340627639681,0.0160363422212768,0.020316074342025,0.0114730598211097,0.00182335331842109,0.00123704493265708,0.00830093726495451,0.0114724478680432,-0.00456864864310824,0.0029851108523391
"1259",-0.00491598804806048,0.00476470863053735,0.00774339094091769,0.00079110445869901,0.00322676566722802,0.00351708159957709,-0.00490460039626495,0.0028357378902979,0.0109751832107272,-0.00148807495388825
"1260",0.0159361874167991,0.0314166312569657,0.0197583959758065,0.0305748357038502,-0.0150098915227197,-0.00634679631820356,0.00616086080452227,0.0248189556502272,0.0258569173676915,0.0298061975373973
"1261",0.00156874237093563,-0.0103447860482367,-0.00107613371275805,-0.00562674497052351,-0.0118896037376056,-0.00314564959670971,-0.0111967840701843,-0.00367841978530026,0.00506675865914263,0.0075978046715317
"1262",0.00266244333115773,-0.0185829552812609,-0.0118537070789172,-0.00437259397330758,-0.0017796789035418,0.000191470706967012,0.0072543714031239,-0.0101541806924524,0.006827847311627,-0.0136445958527361
"1263",-0.00257742255508675,-0.0121304498027494,-0.0109049755661637,-0.0126580483847509,0.00789416723983116,0.00391995887298791,-0.00175672141935257,-0.0059058090929387,-0.00367601726249223,0.00436834231689986
"1264",0.00242770448115648,0.00509153742052315,0.00330786484082957,0.0104656418523008,-0.00176825346786491,0.000190430390057061,-0.00281515987048742,0.00250146727083589,-0.00445290720966107,0.00108748494039279
"1265",0.00867032396069023,0.0146008419225705,0.0120878002733418,0.0217502980458826,-0.00168744930186793,-0.00199956713926652,0.0111166483103398,0.0155956737118539,0.0136741150159743,0.0072410675824528
"1266",0.000542150379377215,-0.00616745899465754,-0.00434340153902912,0.000760482428306508,0.0130155007890431,0.00582022361529466,0.00890059892590767,-0.00061430949860819,0.00649268158404359,-0.00287566377870796
"1267",0.00239928877028994,0.0100472460926062,-0.00436188507683333,0.00405169871086031,-0.00141831248970847,-0.00208704291104933,-0.00657319351782792,0.0129072514091939,0.00444671515559247,-0.014059040274147
"1268",-0.0051731839616721,-0.0184317467224289,0.00219045064284362,-0.00907926433671713,0.00994211330661021,0.00446787915459357,0.0045273398175929,-0.00697814985026324,-0.00698347652501952,-0.00219379185917579
"1269",0.00388075161477675,0.0157972734793712,0,0.0190886778802386,0.0046325766711075,0.000946391320027828,0.00520022199377745,0.00824937730009734,0.00778604193727372,0.00696219963645928
"1270",0.0110561873623554,0.0184857551414892,0.0120219991407855,0.0252246956659283,-0.012104220394993,-0.00311995051263969,0.00638033528146664,0.0139394749145756,0.00685361993769473,0.000363970964420313
"1271",0.0052763174000412,0.0164218706483028,0.00755948299156151,0.00876973465806841,-0.0137535730616226,-0.00597524838008012,0.00633969991109296,0.0197246877076409,-0.00235151600180017,0.00436516390143638
"1272",0.0037273516117291,0.00255109104321161,0.0128617021266892,-0.000724584891686142,-0.0113256792785338,-0.00343448527934753,0.00476755194752543,0.00820666961298255,0.00527233590576648,-0.00724372798843753
"1273",-0.0025766171028726,0.00763351129595891,0.00423261305786959,0.00966657412428784,-0.0063258555053205,-0.00220226975335569,0.00305058641867362,0.00668590664732149,0.00672547018523906,0.0116745244053
"1274",-0.00113982985627337,-0.00280558117970198,-0.0094835990950668,0.00143599421100227,0.00180686451713785,0.00115151509642719,0.00557535674827103,-0.00779676931600581,-0.00704835113879987,0.00180315100471051
"1275",0.0083673863298146,0.00675253207889681,0.0127660461584185,0.0112335537851562,-0.00240424549863694,0.0047916016446059,0.0127686009277732,0.0130968764171717,0.0272205612993197,0.00827933561250238
"1276",-0.00512978695554622,0.00251569031269283,-0.00210095404887267,-0.00401811466168123,0.0132560534893353,0.00534204155648776,0.00580654885094689,-0.00229836602281563,0.00510759530233873,0.00285608377297009
"1277",-0.0004548171613038,0.000557454502880139,0.00526327918843417,0.00522063198869671,0.00314335388617848,0.00303642070409937,0.00247386243425307,0.0051829385646931,0.0101631910046465,0.00356001051713029
"1278",-0.00341349969251337,-0.0153247317994962,-0.00628288436285618,-0.014400241155349,0.0117717369446102,0.00340448878694888,-0.00872001913332132,-0.00773418959027383,-0.00556312951670035,-0.0102873049938557
"1279",-0.00038075942956739,0.00679143206520849,0.00632260858144496,0.00862289683904205,0.0115511033147604,0.00377128791215298,0.00514518520020002,0.00346431372271327,0.00761768141175789,-0.00250900001479271
"1280",0.00875720211993869,0.0207978573737269,0.00628276557974194,0.0220846936939343,-0.011454983241066,-0.00347179158082567,0.00743074632303387,0.0161102929025081,0.00147658143614171,0.00323395006293814
"1281",0.00158530126002554,0.00220306595823283,0.00312187273055997,0.00278835344089257,-0.000419471399055737,0.00141597726976905,0.00213086226016124,-0.00141535186260178,0.00878747946198954,0.00250709217230694
"1282",0.0140185163874254,0.0189558661749092,0.0031119216243265,0.0166818631322894,-0.0214886659827969,-0.00791928199930403,0.0143929288084452,0.0144599369925984,-0.019935714353656,0.0117899484229973
"1283",-0.000668780965979665,-0.00620100680608915,-0.00310226761066446,-0.00843192820911376,0.00995102795471925,0.00275579307854135,-0.00483698967274704,-0.00614884518322967,-0.00274401099226917,0.00494350813762146
"1284",0.00252890738980449,0.00678231922439765,0.0103730916934424,0.00206840104522166,-0.0124013500671702,-0.00644442300837011,-0.000810137910396413,0.00337455611248227,0.0150735979514007,-0.000702731107745658
"1285",0.00296719529622491,0.00323361627290297,0.00410682448898214,0.00711024471247157,0.000773926480035936,0.000476932744866376,0.000648784446100059,0.00532482676417234,-0.00707128474492547,0.00457096435919468
"1286",0.00125749367625527,0.00268610279935566,-0.00306728861869998,-0.000455779826920688,-0.00747680603643874,-0.00228802114185223,-0.00729220324730606,0.00139394942607018,-0.00284864094955495,0.00525029928143272
"1287",-0.00738731300345796,-0.0192876606530892,-0.0123076304650366,-0.0221003337761296,0.0129879193970526,0.00563746795990627,-0.00832523984829647,-0.0153115872343019,-0.00523750136323065,-0.00940102202020787
"1288",0.007442291540531,0.0101065541264962,0.010383981561106,0.0163090728263446,0.001282444987877,-0.000664875325532388,0.0113579204640026,0.00706818494976313,0.00221368913613551,0.00246042320711748
"1289",-0.00125591437187478,-0.0089235089235089,-0.0030830505522883,-0.00825301449791938,0.00529283285201232,0.00209163747837948,-0.00992809405903661,-0.00561505906479343,-0.00232821928028837,-0.000350626340403282
"1290",-0.00465973104768957,-0.00300159691194601,0.0164948594667127,0.00277392537120047,-0.0017834295035829,0.000759258622940573,-0.00493205557131104,0.008469954212732,0.00592392310686707,0.00350749322354549
"1291",0.0110731027256314,0.0139573809003248,0.0101418453607813,0.0108344572487018,-0.00799647311083951,-0.0045506233814433,0.0082603381664319,0.0089583514576641,-0.000654339416725214,0.00454391175146429
"1292",0.00264621720122848,0.0043182878640744,0.00100397078131831,0.00182431109830894,-0.000256948656213507,-0.00104795046658845,0.00163859464203764,0.00721443083543027,-0.00386901190476185,-0.00173971176077381
"1293",0.000439910906924634,0.00134370530903904,-0.00100296383493326,-0.0040972524571673,-0.0110658130605799,-0.00362331028190144,-0.012432488060361,-0.00688709934497111,0.0219300739074966,0.01568487205973
"1294",-0.00322444863180138,-0.0050990578489738,0.0030119692906807,0.00182867127329756,0.0125769973442369,0.00392353686207181,-0.00811657490350237,-0.00693490294372123,0.0112267451473103,0.00926559358588586
"1295",0.00441097641156007,0.00971114525856986,0.00600604786318049,-0.00182533333865698,0,0.00142977658431964,0.0116901536923293,0.00810071441323545,0.000462599740226777,0.00306014184494452
"1296",0.0021954462092495,0.00854923570499344,0.00199024225393507,0.0100569981186751,0.00651057773261043,0.00076113210569595,0.00280608868063537,0.011914800090973,-0.00456599226526433,0.00610175144674652
"1297",0.00167996031185003,-0.00741721216950575,-0.00595844473763918,-0.00995686197650947,0.00885095696175497,0.00332878191688968,-0.00115233383825564,-0.00492919329959496,-0.00307727464616558,-0.00808621224280259
"1298",0.00291637805864631,0.00854061817055407,0.0159840316637869,0.0139430232148705,-0.00329014519362192,0.000474337239811495,-0.00758072688181743,0.00963148859666774,0.0104252069381223,-0.000339669258072273
"1299",-0.0039256130502715,-0.0108496052873783,-0.0176992088182166,-0.000676184218065257,-0.00609414564154342,-0.00397940452940004,-0.00132847645201672,-0.00572386506510203,-0.0530290606654832,-0.0037377712839286
"1300",0.0051815257230956,0.0136436623839418,0.00600604786318049,0.00947413930597052,-0.00941418385797166,-0.00324019191520675,0.00532097459752157,0.00986861182333887,0.0141214200429116,0.0156890517662007
"1301",-0.00304943846279793,-0.0113487751281974,-0.00995025184479759,-0.00245831123725471,0.0093919879710167,0.0040154217544881,-0.000330839746813916,-0.00488587894469106,-0.00162058098781237,-0.0100739096678047
"1302",-0.00407826634832442,-0.004003941409497,-0.00602985052335769,-0.0172487991709466,-0.00793868682648313,-0.00199925407493118,0.00810733076983539,-0.00436459657716448,-0.00414814245877471,-0.00474902210510297
"1303",-0.0146251642433027,-0.0399359964503607,-0.0080893000179334,-0.033508259345744,0.0121323403668563,0.00419749274822112,-0.0134580922464768,-0.0263014546951795,-0.0178086151937923,-0.0163598703524483
"1304",0.00697555185116983,0.0142380734803238,0.0061163372005324,0.0120283662996061,-0.00612112704898615,-0.00189976975547945,0.00432533136901414,0.0123803100598969,0.00571609107036442,0.00450444281824036
"1305",0.00994908908545389,0.0253231536325937,0.0172238511915803,0.0209742298317772,-0.0100074929957978,-0.00295106331668116,-0.0023190182112115,0.0216787898096147,0.0100836885019957,0.00827878144789507
"1306",0.00386781603950337,-0.00697955952038265,0.00398413824371335,-0.000456521280128186,0.00198688582082585,-0.00076358550136435,0.00464890663567052,-0.00516871968716437,0.00665540904317163,0.00273687664164446
"1307",0.0000728068708331087,0.00162189852859096,-0.00992072122176646,-0.0109615692604759,-0.000172640670854318,-0.000287145196488092,0.00694102463673896,0.000547242326691233,-0.00787353023579973,-0.00136470329624794
"1308",0.018025607425791,0.0178135031628575,0.00901819771477808,0.0272457132050588,-0.0175935202680416,-0.00716676872844824,0.0178891023394376,0.0177643773340344,-0.0167807831982463,0.00444138199630006
"1309",-0.00107080293416262,-0.00689435375724667,-0.0109236886218586,-0.0157339729339958,-0.0251956880858202,-0.0114546804338819,-0.00241857090709896,-0.00939879888135564,-0.0168206774463214,-0.00680273323384251
"1310",0.00578919669838163,0.00961281027826755,0.00803213640426526,0.00799263534092987,0.00153168518057112,-0.000292573833753362,-0.000646360471140861,0.009216643676208,0.00946289987942417,0.000684922163946666
"1311",0.00138503976134308,0.00872768686346315,0.00597624973529531,-0.0011325548789618,0.00197785367547731,-0.000291353956402896,0.00598414567439742,0.00637937694001067,0.00136578716953339,0.0123204071609913
"1312",0.00392000886614152,0.00471948539726963,0.00297021874301184,-0.00385597609196009,-0.0119354259576846,-0.00613848723071353,0.0059483969913241,-0.00134282171204159,0.00179784869563826,-0.00169030813224702
"1313",-0.00291091567169599,-0.0117431751769635,-0.00987178217331175,-0.0173040634105102,0.0039960122488647,0.00049051391830246,-0.00239731129209275,-0.00995158596000634,-0.00903515710217606,-0.0121910687751201
"1314",-0.00163767979038254,-0.00580942994098665,-0.00498501811302132,0.00185344840426627,0.011308328028532,0.00509454519616193,-0.00224285731284235,-0.00353163525869626,0.000499606554061893,-0.00239976354492633
"1315",-0.00720382457959412,-0.011420950456558,0.00100193040466778,-0.0152637138837692,0.00322024140051447,0.00126743623858006,-0.0118815139323681,-0.0109053543489495,-0.00399475670705129,-0.00790370781297056
"1316",0.00323283015856712,0.00698532089438597,0,0.00751531264627725,0.00945143425702244,0.003699768676938,0.00406212064991829,0.00303195916485222,0.0122829599173986,0.00969855199605174
"1317",0.0140353565933733,0.0170758310782111,0.00700708895954683,0.0174826083987241,-0.00512308959118413,-0.00116378782864435,0.0103337338566905,0.0129157692033499,0.0177675665063304,0.0044597718600301
"1318",-0.00310687835597034,-0.0115422959647333,0.00795229407247633,-0.00526921146169612,0.00719198398501164,0.00553546313085462,-0.000485048641219232,-0.00189901952320193,-0.00705589441809829,-0.00409837491775156
"1319",-0.00495890188087655,-0.0111467704919681,0.0019723535448064,-0.0168126403611232,-0.00141067059251088,-0.00173852231321836,-0.00226284416491651,-0.00679548338608327,-0.0105979536082469,-0.00960224010502808
"1320",-0.00170889661567153,-0.00778303269008052,-0.000984179686273512,-0.00117102311228512,0.00750352379203312,0.00416042842027187,0.000972054773094255,-0.00191531691132452,-0.00142403570751148,-0.0138504051469359
"1321",0.00413646014301605,0.0102786603360474,0.00295589479626401,0.00727001674528394,-0.0169107767096219,-0.00491418721008685,0.00841707230740241,0.00959679982476702,0.00520830856403953,0.0112359826673936
"1322",0.00731489596847457,0.0152609565133073,0.000981827964540827,0.0137369569146719,0.0055401229019536,0.0023961283668279,0.00642037731267631,0.0103202907782867,0.00505802507580877,0.0128472255229006
"1323",-0.00408925071169619,-0.020833130241711,-0.0127573945941051,-0.00574198543754867,-0.0173284003478921,-0.00735380937949048,-0.00462528980260168,-0.0129030889534346,-0.0187185648862335,-0.00445657267375199
"1324",-0.00991110804519513,-0.0258552689559963,-0.0228628066966687,-0.0180178963725313,0.0137455185116302,0.00506888629287983,-0.0100943874085713,-0.0152502839994878,-0.0167614736178715,-0.0154959387610798
"1325",-0.000500469299067885,-0.0091236253856225,0,0.00541040526272418,0.0072258259476079,0.00446116175810984,-0.00437031224624473,-0.00359545476145628,0.00699695280848123,0.0038475546290011
"1326",-0.0112308043620832,-0.00446418523737035,-0.0061036905276256,-0.0147400475654865,0.0233809436704899,0.0102346034835701,-0.00959222631567447,-0.00499614279578853,0.00669570471474579,-0.00452973397957102
"1327",-0.0167848892084438,-0.0252243080852308,-0.0122826970358146,-0.0194728013399279,0.0113375769201478,0.00468311594177906,-0.0193693790726244,-0.0108781976195985,0.0108553118797552,-0.0133005924675427
"1328",0.00809411204075516,0.0169639268328183,0.0134715136150008,0.0108983693632969,-0.0119804421882446,-0.00389991076162077,0.0118846598428499,0.0118443535208888,-0.000186213525032453,0.0024831161464689
"1329",0.0130657747847533,0.0197907790473342,0.00511259232487116,0.0256346799699372,-0.00415668764789889,-0.0020055822589583,0.0142266529599688,0.0139355777469419,0.0101197611545394,0.0130927143080344
"1330",-0.0118885397249796,-0.0263376411996569,-0.0111901618088022,-0.0151833547890955,0.0161764423646942,0.0060283147970801,-0.0052193109535672,-0.00769675817123416,-0.011370565667558,-0.0101291689588564
"1331",-0.000656356454987184,0.0105350435304219,0.00205737429440145,-0.00498082074390671,-0.00145533009479659,-0.000285575947685301,0.011641323832565,0.00332397916059901,-0.00242461290302975,-0.00988007454080853
"1332",0.0148125505581382,0.0208511069798401,0.00616029496647896,0.0114421358154058,-0.000599658427548833,-0.00104614886263132,0.00858992824453608,0.0124240360459011,-0.00130878094751663,0.00463293958054045
"1333",-0.0033796017364337,-0.00800426385435349,-0.00204089794416418,-0.00471366476542112,0.00291609408232896,0.00199996790564905,-0.00530296976829436,0.00245414023793811,-0.00586584711388449,-0.00957784323772171
"1334",-0.00642077129957053,-0.00528693460894625,-0.0061347802193088,-0.00449910321548197,0.000940843647144085,0.00114060354514489,-0.000484732868428983,-0.00435256650663762,0.000753217007761098,0.000358161290763714
"1335",0.00167008361232535,0.0125875148132877,0.00205737429440145,0.00689823205459028,0.000170605570384508,0.0000951638765260832,0.0105060477358532,0.00928984569977431,0.000689958005580582,0.00393840047884164
"1336",-0.00840906436449851,-0.0223755753006758,-0.0112933305971585,-0.0191355533462609,0.00726053206286803,0.00199343495803439,-0.00927721221427358,-0.0143474329231922,-0.00294588203974666,-0.00178321596697351
"1337",0.00380148767320909,0.00734667204270645,0.00623033592831779,0.0021677378288214,-0.00703862107838005,-0.00255840224745696,0.0127545062560026,0.0120842789233824,0.00144587910906413,0
"1338",0.013691760118048,0.0165496541470023,0.00515984322393015,0.00913248214632767,-0.00512432507296423,-0.001234623465596,0.010999444840446,0.010854880824958,0.00200873819192582,0.00571639657127987
"1339",0.00696867357320885,0.0066227008726909,0.00513355972773066,0.00619186979810071,0.00600864775653021,0.00332851402223411,0.00425738324519531,0.00375872403197142,0.00883350485006607,0.00213140957556313
"1340",0.00164114344063737,0.00520818715348192,-0.00306435818446671,0.00142024517741746,0.00085390294508958,0.00104371521895996,0.00486730587994466,0.00401167278015757,0.00217354531561553,0.00319035098056442
"1341",-0.00370388151839296,-0.00627189261221206,-0.00204926237770342,-0.00212717758902492,0.000255661752853298,0.000851724251571317,-0.00140633646115407,-0.0037293620130171,0.00309827726179579,0.00388694552119162
"1342",0.0062199597313255,0.00768371518461985,-0.0102665953584101,0.00663142931494987,-0.00518634994809586,-0.00181949692206418,0.00876237826339032,0.00267355719597395,-0.00345934014518967,0
"1343",-0.00298430479014788,-0.0106207592448013,-0.00518692828762368,-0.00188214830567857,0.00704249970042459,0.00189838404920217,-0.00155131731176716,-0.00239990331815743,-0.00452523536029847,-0.0130235865097412
"1344",-0.00762530584787435,-0.0090834423099786,-0.00834194245807418,-0.00754346341545686,-0.0002557684276141,-0.0000946584414326379,-0.00341755307609259,-0.00908837443434851,-0.0100877703490323,-0.0110556673761554
"1345",-0.01615813224316,-0.0172224263141999,-0.00736063863969971,-0.017577174661878,0.00784889649385123,0.00398076482564025,-0.00763835471815877,-0.012948499535044,0.00314524751119549,-0.017670375073744
"1346",0.000730073787724717,0.00819674544411231,0.0042372467644598,0.00362681492579564,0.000168706606664237,-0.000283610830367875,0.0056550125769923,0.008198685224452,-0.00244559476738193,-0.00220261312828607
"1347",-0.00401176072440168,-0.0134567390961072,-0.00843894592525607,-0.0158998535536409,0.0053321836543101,0.00226631651311116,-0.000937299617321252,-0.0103006686917689,-0.0193613399627692,-0.00367920130409782
"1348",-0.00593173909213995,-0.0147769629821647,-0.00851040579899298,-0.012974483048442,0.000673779896261273,0.000847978439536767,-0.00234508179475645,-0.0106819626231863,-0.00980768589743597,-0.00775473278825167
"1349",0.00206277523301424,0.00519187970960644,0.00429143816809052,0.00421640099469545,-0.00294526851158161,-0.00141227856578552,-0.000940300479815304,-0.000276960878379695,0.00194214409307869,0.000372080552337062
"1350",-0.00301440948795484,-0.00487794120648877,-0.010683523668543,-0.0128426287987381,0.00826902807783036,0.00329955374173463,0.00423526127838336,-0.00498465198157827,-0.00781809115931786,-0.0074404513480204
"1351",-0.0110610202980634,-0.0204728873617209,-0.0107989857845252,-0.0227669734861317,0.0139748835489482,0.00441523015989786,-0.0121835799710409,-0.0125243124105806,-0.0145219850810365,-0.0131184545155544
"1352",-0.00574174385333626,-0.0156019594506337,-0.0131007105903591,-0.00870473395400018,0.00404420134593275,0.000281113784746045,-0.0049019403780779,-0.00930113876704308,-0.0105068193946103,0.00189894864774565
"1353",-0.00382452313896431,-0.00687807899270176,-0.0110617943502787,-0.0142046259009562,0.00287658000496438,0.000747554040916087,-0.0122358307793132,-0.00825030652236147,-0.0018698944213339,-0.0011372096858524
"1354",-0.014831056042912,-0.0165613401065168,0.0089486811943067,-0.0136232144509609,0.0177035990775352,0.00373763753562839,-0.0276704746990554,-0.0117615060852646,0.0223470884756483,-0.00227693068930646
"1355",-0.00855895077693458,-0.00275562422834985,-0.0144125503521981,-0.00956175397065728,0.000241888644155974,-0.000651145360915706,-0.0102581744298914,-0.00725662154666429,0.0114528793562916,-0.000760813374248825
"1356",0.0171883904314187,0.0239484975494237,0.010123309457468,0.023867068097517,-0.00209360962528693,-0.00260843197606475,0.0205615340118657,0.0236839186567812,0.000646981546807091,0.0133231960579028
"1357",0.00174265531466289,-0.00329837850990267,-0.00111309381846691,-0.0104764505845661,-0.0111341350985775,-0.00214806391720246,0.00212961601768935,-0.00628397537980041,-0.0166181189764546,-0.0142750178179645
"1358",0.000529670840551999,-0.0105293280307589,-0.00780375375636477,-0.00688229851231248,0.00693509443252593,0.00262030723866213,0.00424950365411148,-0.00546093508726975,-0.003024769818191,-0.0110518353072266
"1359",0.00196569671129598,-0.00638513371548355,-0.00449468849517021,-0.0050636677956738,-0.00380832119563679,-0.0021464872984247,0.00309266997694935,-0.000867559826956521,-0.00138498223799577,0.000385351197087491
"1360",-0.00324449326236353,-0.00152988765638218,-0.00564321528067357,-0.0048219061492506,0.00374151668039047,0.00289958425634862,-0.00292074819724564,0,0.00838774827586697,0.00346682482868865
"1361",0.0121117274077596,0.00950047561552636,0.012485860502307,0.0282635278036116,-0.00307925853634017,-0.000839250190217244,0.0136696066990811,0.0138851665676218,-0.0108723413420644,-0.00422251234308701
"1362",-0.0145099174472471,-0.0258045756486026,-0.0134529437399317,-0.0172774115122138,0.0253615547248338,0.00952274148181065,-0.0232781341913977,-0.0199712471827835,0.00589325901487858,-0.0185043039401039
"1363",-0.00220111584753857,0.00124663432088945,0.0102273272562641,0.00426219469363875,0.0115743199169493,0.00388426946179066,0.00624567936413678,0.00378424444983616,-0.00190908427597691,-0.00864096828130689
"1364",-0.0251766722562305,-0.0211641431203992,-0.0269967785366355,-0.0267903376331318,0.0237402014110479,0.00858997028705999,-0.0253184020318392,-0.0179813425170152,0.0387811976909775,-0.0206023441985491
"1365",-0.000468200518593642,0.00699524913418226,0.0115607965464521,0.00436080666081362,-0.00790091184935682,-0.00576295041738184,-0.00703862369897512,0.00383945835388255,-0.00114281269841265,0.00566352009082416
"1366",0.00757246509894727,0.0031574357857429,0.0125712831486959,0.00271360172024693,-0.0133769582786138,-0.00331266301139854,0.0197468540118362,0.0061783213547264,-0.00114421556058042,-0.00362030687199211
"1367",0.0224682128837408,0.0336794815837116,0.0158013484769939,0.029228656216727,-0.0199842114251529,-0.00655470393045698,0.0213506492311568,0.0362571072869038,0.00044551355762712,0.0185708895967318
"1368",0.000606097106397474,0.00182716848995401,-0.00666646163817064,0.00604791734863563,0.00151931082413559,0.00241646019864894,-0.00486164593552263,-0.00423257848789793,-0.0172381329389546,-0.00673799981177947
"1369",0.00795147755599457,0,-0.00894874463830775,-0.00862525052444796,-0.000239181574910985,0.00074109201463135,0.0125387547801934,-0.00510047602802599,0.00148864724919084,0.0031922947283809
"1370",-0.0126974244539807,-0.0112462681363305,-0.0045143737722364,-0.0145002577141462,0.00455211658883226,0.00268690270845573,-0.0196205286374211,-0.015095248312049,0.00407164102815605,-0.0182974890606896
"1371",0.0114913120756084,0.0190595215836558,0.0113377413974922,0.0208666605454313,-0.00914269872053086,-0.00535867655892219,0.00935031886285587,0.0118562109314444,0.00708036813156299,0.00486217012124057
"1372",-0.00639499137092681,-0.00904987050920769,-0.00560538262726251,-0.00366879961400224,0.00986905889919476,0.00529433623064279,-0.00471324061517497,-0.00600174921678587,0.00421825367807882,-0.00766118603546284
"1373",0.0106002335643784,0.00700165174665401,0.00789179765816006,0.0071015651348687,-0.00127146158086444,-0.00267921162740137,0.0135532379913388,0.011213518364847,0.00400970608483031,0.0117837915331112
"1374",0.010227554452708,0.0157193129592765,0.0145413333384934,0.0182814066227075,0.00556892387400709,0.00463189505477857,0.00628353741616117,0.0120371367792191,0.000570497622820909,-0.00160644505840102
"1375",0.00193828235965432,-0.00922620706164989,0.00220537871899129,0.00205195096251232,0.00537969259920157,-0.000276721574093863,0.00784479173446284,0.000855674030864506,0.000570178676385646,0.000804494238004771
"1376",0.00967246457235493,0.023130189836249,0.00550030036382165,0.0161247594875984,-0.0130625697118006,-0.00341274212644982,0.00466377173952437,0.0170985074790255,-0.00487550835261552,0.00844052334810597
"1377",-0.00162126786648054,0.00703774436524318,0.00875277447287925,-0.00327435229046324,0.00494332169447609,-0.00203647153836795,-0.00127636589375379,0.00196165230000989,-0.00757192014324448,-0.0163411536663084
"1378",-0.0224387118095651,-0.0275945539306232,-0.0144548389171494,-0.0366220805818028,0.00531549205039372,0.00213353800312532,-0.0156522854387714,-0.0209731077196352,-0.0253253636896495,-0.0214749183216139
"1379",0.00770148081128275,0.0111042254999525,0.00666700061124326,0.00318541991386323,-0.0133372680529092,-0.00434996372525542,0.00081129607158914,0.00942585690894071,0.00407837773770869,0.00993788052228783
"1380",-0.0160345538783295,-0.0265405595701065,-0.0154527701620444,-0.0185234906933806,0.0145577329640842,0.00548408863164052,-0.00551256020272284,-0.0116015301925666,0.00733750004807066,0.0102500893865118
"1381",0.0050257544284229,0.00626753714331851,0.0112108294768711,0.00862767929779129,-0.00394178296583025,-0.00221882655222094,0.00440209215883569,0.00973380237703614,-0.00741415216617314,0.00689934024072114
"1382",0.00901674449582557,0.0084087746584518,0.00776069645006561,0.00641543296342362,0.00158280794044874,0.00138953341528425,0.0063299734012543,0.0110571896152669,0.00137601236325557,0.00564301657149979
"1383",-0.00285360525269862,-0.00154421688393624,0.014301302392695,-0.00478080942116232,0.00244992905117813,0.0032383788338548,0.00838707524348847,0.00168289076484562,-0.0116469212635357,-0.0108217008893704
"1384",0.0249266360563531,0.0423755687483474,0.0206073625167946,0.0443020698938861,-0.0130075692597558,-0.00461105179269228,0.0227126561764064,0.0296751689788228,0.0274081358343303,0.0433548923793641
"1385",0.00301262298268568,0.00919873054601927,-0.00318821209263942,0,0.0103175218466918,0.00463954765149222,0.0106352866263599,0.0103318964143853,-0.000644410069663981,-0.00194172110753565
"1386",0.00659258782972572,0.00793886465006532,0.0127931580728333,0.0199336954493066,-0.00768509946474538,-0.00249341323488661,0.00557104508706852,0.00430564072935535,0.0152815208016381,0.0280155820911756
"1387",-0.00451175506974522,-0.0239205878540124,-0.0126315605223641,-0.0105238531041365,0.00510986603831354,0.00268487196029055,-0.00461710587067177,-0.00911060279757225,-0.0113045466840351,0.00378503751243242
"1388",-0.00950366181868567,-0.0128510228128618,-0.00426407658837935,-0.0182323870145652,0.00929413883510399,0.00350928366334946,0.00139139288567525,-0.00432643728942272,-0.0126540730252988,-0.023001542465737
"1389",-0.00125463963770434,-0.000605568531430678,-0.00535371043379596,-0.00361130209659422,0.00881417770635795,0.00276019569632413,0.00200730170336261,-0.000815098654200819,0.00214680882813312,0.0177537984865639
"1390",-0.00872015260636338,-0.0042413238337734,-0.0107642979607504,-0.0111310505309794,0.00202884278508764,0.000459108198425984,-0.0118645012565484,-0.0103286412550253,-0.0122695344448635,-0.0128934580304473
"1391",0.000148846071287068,0.00365098559631694,0.00217659142597859,0.00523550809382511,0.00124563405599987,-0.000917550697881686,0.00155933819713883,0.0107110296875805,0.00552094007969539,0.0111409573662571
"1392",-0.00484482016187215,-0.010306436106676,-0.0152010057799163,-0.0166664547702504,0.00707620756684868,0.00229569102181792,0.00435939874862279,-0.00624979714408214,-0.00261460871251018,0.00227960414753747
"1393",0.0167775766206038,0.0159267098827598,0.00992302401152001,0.0193325300154563,-0.00262535390182472,-0.000824420053331165,0.0108511305958692,0.0150394798913043,0.0101579595034524,0.0121305097542026
"1394",-0.00235726487658972,0.000602938215416904,-0.00436719305748223,-0.00233838962562882,0.00464504791081599,0.00219988873732957,0.00383343559525318,0,0.000454184510537026,0.012359496595415
"1395",0.00686709132876984,0.0042180242998735,-0.00438597950133768,0.0132811874123728,-0.00785992558009407,-0.00256112386589702,0.00840212932917384,0.00942931813235459,-0.00479868988009313,0.00110978658825989
"1396",0.00740681658627573,0.00690085679541297,0.00330405313311677,-0.0025699876669133,0.000543559942194571,0.00100902190980912,-0.0077261467185249,0.00400287225516593,-0.00273667816031353,0.00886924934503464
"1397",0.00262087725885984,0.00953508736428077,0.00768402762864495,0.00927616408397958,-0.00256151667350246,-0.00146618592204739,-0.00839683641550082,0.00318990545196018,0.00215617114362288,0.0120879356194799
"1398",-0.00914841253302245,-0.0242030009194759,-0.0239651238801355,-0.0148073616400825,0.0122188902861524,0.00394560990847248,-0.00338720468292908,-0.0116586646127462,0.00189068320867491,0
"1399",-0.0101122828153909,-0.022988519914049,-0.0133929609867391,-0.0261725927976761,0.00561277946488237,0.00164474474550125,-0.00602503243833441,-0.0131368060232953,-0.00416476220686868,-0.0209916867428366
"1400",-0.00858706556297295,-0.014551168722522,-0.00904992960961082,-0.00425763898236642,0.00787534303099591,0.00191640309022345,-0.00404102193767331,-0.00869336549230293,0.00320201923284325,-0.0059150056241617
"1401",0.000224413245655475,0.00691168773141393,0,0.00481047774018739,0.00257893099894102,0.0005463502855938,-0.000156134047395007,0.0112362322794795,0.0140046504949283,0.00743779921520837
"1402",0.0164969752562591,0.039001532955854,0.0148404084932059,0.0226063026798382,-0.00915571758241562,-0.00309508143940618,0.00811616533119142,0.0181567983994437,0.00706626847904257,0.00184567420582926
"1403",0.0184332665999447,0.0252252896308165,0.0179977431019347,0.0280881839021998,-0.0188620249544126,-0.00721218726737272,0.0113020060149582,0.0159703557223849,0.00491158372363132,0.0103168479898337
"1404",0,0.000292921742659713,-0.00552501877991773,-0.00581835466358038,0.00747239807680522,0.00321889230229422,0.00275562188802891,-0.00314398047599751,-0.000698235399820168,0.00583515216558039
"1405",-0.00699444011399852,-0.00732060985955085,-0.00111091188872348,-0.00458002932519108,0.00200830180246347,0.0017412536393473,-0.00106849596260239,-0.00210238718666944,-0.00597083174614632,-0.0119652153326775
"1406",-0.000871358929212196,0.00147497755845039,-0.00333703580461586,0.00178933100786272,-0.00499901544389236,-0.00364697323657004,-0.00290406324899295,0.00237020811570932,-0.0086267873785294,0.00146794543273732
"1407",-0.00690493027736772,-0.0191459584690391,-0.00446439347680483,-0.0117375144578268,0.0056682916667834,0.00239136081218638,0.00107289634318009,-0.00236460351327161,-0.00651021017474662,-0.00842810650609738
"1408",0.0198333914289337,0.0441441641539726,0.0112108294768711,0.03098363004042,-0.0161372879264327,-0.00523057774482527,0.00734998500516326,0.0265999813709239,0.00921298873635923,0.0169993723911357
"1409",0.00193770924393943,0.00603958039920172,0.0099776868493977,0.00626121259229673,0.000391994865878154,0.000645687644220683,-0.00288809135276169,-0.00307841797263331,0.00482160067846471,0.00581391130596076
"1410",0.0050135033486447,0.00857634695033704,0.0120748212746327,0.00273738760263686,-0.0128655216410212,-0.00525444247299922,-0.0103659181400872,0.0038598469460116,-0.000127984642457113,0.00758667603917651
"1411",0.00121146170529118,0.000283596618301907,-0.00216938686191614,0.00198529434522365,-0.00532421517857529,-0.00139033510807585,-0.00600750079087131,-0.00589580892404773,0.00127973509905122,0.00286844636302375
"1412",0.000854240735612466,-0.00113360999869283,0.00217410333312351,0.0042114078973805,-0.000719613026230803,-0.00074243069037172,-0.00294432027845992,-0.00567327248365324,0.00325926005263955,0.00822316790061595
"1413",0.00163584701576558,0.000567465778748666,0.00108464773335926,0.00468676977792315,0.0050371291436333,0.0028793557851674,0.00217605525163522,0.00207485325255097,0.00121019169341396,-0.00531922193021361
"1414",-0.000497197239003766,-0.00255179765900493,-0.00216682336640328,-0.00883908932222821,-0.00167011547034024,-0.000648209528922195,-0.000310577437989235,-0.000776395827119969,-0.00757086176992006,-0.00784314027661215
"1415",0.000141959552837356,0.00454812729238929,-0.0010860388260252,-0.000247229342661193,-0.0135472010359691,-0.00491096216271913,-0.000465168342092648,0.000776999085968066,-0.00551317374468951,0.00107795869947758
"1416",0.00113650573072088,-0.00226390750050254,-0.00543472403506051,-0.00148683255435178,-0.0140562263978158,-0.0050286143642243,0.00279385090872064,0.000776434660503034,0.00322310309988061,0.00861456835818042
"1417",0.00737853831334756,0.0116279990029442,0.0131148268680399,0.00918106207228031,-0.00852075907937466,-0.0024331376340988,0.00727435134669241,0.00517193062567833,0.0059756664532653,0.00391453712345635
"1418",0.00133801858225557,0.000841106885306919,0.00755149149820133,-0.00491754223549656,0.00487559912086932,0.0012197422509419,-0.000460818087256398,-0.00154360353794269,0.00102199158178307,0.00141799052216385
"1419",0.0000704638690198767,-0.00224080154889827,-0.00214151424716424,-0.000494225092292133,0.00205589093890879,0.000561921215973316,-0.000768723623107093,-0.00206121680921678,0.00344559722150595,0.00460174330616092
"1420",-0.00302451037334306,0.00842211155264549,0,-0.00148332116548333,0.00443153611907698,0.000842944536361356,0,0.00180728992443613,0.00998351169984457,0.00916132853008333
"1421",0.000423609644229161,-0.00250544909827033,-0.0010729797408694,0.000495320522999831,0.0165044084542907,0.00776686687145833,-0.000923014982832648,0.00180410686655064,0.0107661712426346,0.00523746664346136
"1422",-0.00817944639748758,-0.00586100735454365,0,-0.00915606924300294,0.00417989451222467,0.00176389277894984,-0.00261800598861783,-0.00565975096045745,0.00840915696314992,-0.00486276892515303
"1423",0.00604295681993694,-0.00364958860579034,-0.00107416243358638,0.000249707543371391,-0.000960433761349799,-0.000463262876595927,0.00385980543025322,0.00129378747518993,0.000494175060190116,-0.00453753155768599
"1424",0.000211899727994291,0.00338093405226769,-0.00322580148273177,-0.0102371864436103,0.00584889173002634,0.00259643317101643,0.00215335865132937,-0.00310111657799828,-0.0037661295069078,-0.00455828677532077
"1425",-0.000988910426054312,0.000561971729843513,-0.0086301677809919,-0.00201808551968674,0.00238982383751885,0.000369492426651297,0.00398994405698661,0.000518609662490732,0.00173523796643993,0.00070453633450196
"1426",0.000777824789085724,-0.00336823846738832,0.00326465790504038,-0.00480299095426884,-0.00437067912617706,-0.000646859389730081,0.000305952934962272,0.00259081013634299,-0.00649593545221427,0.00175991964506861
"1427",-0.00720792491021938,-0.0121089583710829,-0.0184382193754041,-0.0116841781229238,0.00518776575931423,0.0018504144308662,-0.00106969806013724,-0.0108528805340987,-0.000435842840422085,0.0010540966616186
"1428",0.00476896138608707,0.00940707891681702,0.00110514652774274,0.00950928391907224,0.0141337195517881,0.0064638477927248,0.00397724806523736,0.00783681598373964,0.0230500679529013,0.0105300477460186
"1429",-0.000920722931040951,-0.000565006129355838,-0.0132451961353797,-0.00560075601580812,-0.00100421376232052,-0.00228788641233746,0.00502841656628861,-0.00596171638562271,0.00158321153584695,0.000347338084005111
"1430",-0.000851035658953614,0.000565325541751927,-0.0123042731220868,-0.00512032580414223,-0.00471266606023213,-0.000368362026003544,-0.000606494475387631,0.00286852100163659,-0.00103354817688583,-0.00486111622344032
"1431",0.0202966159435662,0.0293700668100656,0.0135898538829304,0.0221306659773308,-0.0166511579256524,-0.00681717676624449,0.00788830867873913,0.017680797959259,0.00352991909841038,-0.000348877680432791
"1432",0.00389484345420832,0.0145405662438334,0.0134079911592158,0.0231621750609929,-0.00465441663959976,0.00129840212613397,0.00180645827074621,0.0107305321013311,0.0215295228426802,0.0111692034417417
"1433",-0.00568098368094239,-0.00919434471770775,0,-0.0127950568637192,0.00241906724891372,0.000463829717175734,-0.00646072345279991,-0.0123861337659207,-0.00682741027276867,0.00138079096165633
"1434",0.00278712054964436,0.0136462928451795,0.00441003331665257,0.0119638193076583,-0.00627361245327607,-0.00185208493320832,0.00393155976401904,0.0104940127182953,0.00364636873408197,0.00206822407648244
"1435",0.00333558969459991,0.0037696523206705,0.0109771999454502,0.00443349335475829,-0.0124648377174081,-0.0049166445979123,0.00376576095343095,0.00531917481336985,0.000119142350892609,0.00515995919531664
"1436",0.0152364858779614,0.0160944503816272,0.0162863736468242,0.026974128977066,-0.00393379838631991,0.0028898866004794,0.0121548812915082,0.0191481921151722,0.0201881850903787,0.00684463933566049
"1437",0.00443394235460315,0.011615575566891,0.0106838856587941,0.0116999208340451,-0.026577956032542,-0.00938847933215503,0.00518910617049695,0.00321408480119567,0.00286034093585119,0.0105370807807292
"1438",-0.0033955733702995,-0.00443644784117492,-0.0095137274768935,-0.0108568828963128,0.0120039542147974,0.00206469672021958,-0.00471998743186242,-0.00936424619973841,-0.00814906272149485,-0.02758157108499
"1439",-0.000818101957051232,-0.00786367926625975,0.00213465826896719,0.000477664959672497,0.00501145583569951,0.00252847768034359,-0.00859496287273953,-0.00273643649683875,0.00774652022581646,-0.00726389441688557
"1440",0.0005456259358676,0.00660498939033194,0.00212978216083837,0,0.0065658171049392,0.00233503943504454,-0.0046338534449103,0.000499076050558989,0.000116491962983467,-0.0146341610358031
"1441",0.0000683561691181556,-0.00839878984105313,-0.0106269955429268,-0.00596244821407399,0.00247677960915071,0.000558713939044164,-0.0117134208805448,-0.00299172805206593,-0.0015721671837613,0.005657667601356
"1442",-0.000417776642485101,0.00158800100323697,0.00537038978009718,0.00239907603438771,0.00115322053434941,0.00214253057637359,-0.0003037573033291,-0.00317912444737922,0.00285767771121659,0.0066807125953503
"1443",-0.00150838703797995,-0.00369991776292711,-0.00213636900395364,-0.000957457589125355,0.00781567841983888,0.00223046380132752,-0.00106430918089073,0.000759466759175931,-0.00529195140123473,-0.0104784481678606
"1444",-0.0106419766560696,-0.00822257580203967,0,-0.0148537444880531,0.00987754450369471,0.0037090986862458,-0.0146784646387866,-0.00758739953052301,-0.00163694238578882,0.0010589336079363
"1445",-0.00562141175432473,-0.0131049700395695,-0.0107068795419665,-0.00462046238611535,0.0107510860111584,0.00415724277681773,-0.000933989573961513,0.003312669152574,-0.00562163130241533,-0.00705219856480976
"1446",0.00942191452946983,0.012195009321625,0.0119046927829405,0.0158805275572296,-0.00711828604134979,-0.00211577700493415,0.00545305194657342,0.00990610144724591,0.0148989931676462,0.0124289901219379
"1447",-0.00463216489206586,-0.0222220363557285,-0.0192513984914844,-0.00601244101019549,0.000564373041848087,0,-0.00232413510489304,-0.0128267643197265,-0.00261110021146815,0.00596284678055925
"1448",0.00263930249317901,0.00930988342951045,-0.00327141045483359,0.00992005378515604,0.00371044279368182,0.00185552692786728,-0.00714530786197765,0.000764270255662725,0.00232703474505236,0.0013946092478001
"1449",0.00103898420569437,0.00623967422620186,-0.00437628913803645,0.00143767552585006,-0.00136621296445805,-0.000644928010086199,0.00844815460873316,0.00229102191564712,-0.00110271639514203,-0.00522287761086537
"1450",0.00408334691462464,-0.00269617181753401,-0.00439549436054276,-0.00669862949893318,0.000322051765638154,0.00101386166057194,0.00294787268174601,0.00101613535607448,0.00180126664260527,-0.0171508047357199
"1451",0.00716785956779953,0.0121654735127235,0.0121409595774455,0.0103563847329904,-0.0124710629128673,-0.00396064434042531,-0.00371234606913018,0.00888094185216026,0.00696013556150743,0.0217237170535389
"1452",0.0000682030380554366,0.00213692549205846,0,0,-0.0129534442483632,-0.00453177082463962,0.00434709994551397,-0.000754616762860927,-0.00570247102296839,-0.00522833851815707
"1453",-0.00342101680013718,-0.00799614432709117,-0.00545262643871236,-0.00882005940818342,0.00841874631529005,0.00325183917092486,-0.00417391907052667,-0.00402673871298431,-0.00330200449837803,-0.00280311720481063
"1454",-0.00988783682238925,-0.0163887503014339,-0.0164471613374949,-0.00745533744789451,-0.00180090656001231,-0.00203750358227306,-0.00434634449491278,-0.00657091110109187,-0.00616098797743125,0.00737878512213519
"1455",-0.00637992203402371,-0.00273152165466517,-0.00780373644183474,-0.00605760248081522,0.00705209343841218,0.00241258121276422,0.00124729508411181,-0.000254166160957414,-0.000877296892294877,-0.00174399536590708
"1456",0.000558704185149361,0.00986018191029481,0.00561772646302994,0.00926365190811218,0.006921651765879,0.000925841883249401,0.000155638367153488,0.00610691240542494,0.0028097109063383,0.0115304929006563
"1457",-0.00327899400062193,-0.000270964773239957,0.0011175575162059,-0.00314004297867065,0.00250663910683468,0.0000923673577810646,-0.00435928299154964,0.0012642280667281,-0.00735471018279843,-0.0138169849865292
"1458",0.0083278961660016,0.009223841487499,0.00669638644608028,0.00581533714859672,-0.00225869235472709,0.000277460420216702,0.00672397309284678,0.0101037968173685,-0.0100552276849962,-0.00490368285955811
"1459",0.0101336026248056,0.0185485700841777,0.0144123215999725,0.0103588792196971,-0.0138246196391965,-0.00471475110746811,0.00465995587679169,0.00975258952106217,0.00635575860923931,0.000704040312520915
"1460",0.00453469260323036,0.0102928546184431,0.00546442165878713,0.00786855354947869,-0.00926407926142925,-0.00631634938997061,0.0015460460799992,0.00990542113177373,0.000708269398043582,0.000351663888966014
"1461",-0.0025989829863754,-0.00548585873404117,0.00652160777947275,-0.00283918650693982,-0.00612293515400741,-0.00177593703954237,0.00941643256140545,-0.00662084039373845,-0.00442373499449178,-0.000351540264949435
"1462",-0.0166643422888428,-0.013396387238898,-0.012958703974295,-0.0154213007679753,0.0135705985263379,0.00421414152519417,-0.00932859051790069,-0.00987371133169024,-0.0107825823536826,-0.0151249139891453
"1463",0.000139552763020578,0.00559098596475827,0.0142231932353092,0.00963892286693135,-0.00640694323774005,-0.00335725168493339,-0.00355044121872738,0.00772815281411399,0.00365335686857904,-0.00464283041474622
"1464",-0.0138763524184208,-0.0238284818497299,-0.0204964250118485,-0.0205251170385472,0.0143022661356238,0.00477157026715402,-0.0100701081494502,-0.0113802148586331,-0.0128297468333961,-0.0121995151716672
"1465",-0.0028283901412689,-0.00135582855575545,0.00220292894394114,0.000974606987582449,-0.00986192350335635,-0.00214163414663759,0.000626267694406879,0.00400400765503783,-0.00344551788743641,-0.00290588105193434
"1466",0.00290714444888107,0.00624662028871392,0.00769209969754869,0.0109541972064777,-0.00510414838582951,-0.00363917586476059,-0.00437913653853172,0.00822518785289028,0.00703629135608219,0.00255005608008707
"1467",-0.000565448513878852,-0.00026994820593762,-0.00545262643871236,-0.00770528873184073,0.0147278420069885,0.0063690862529695,-0.00581210501707663,-0.000494410517579147,-0.000542169605055598,0.00218020271517072
"1468",0,0.00242982318351803,-0.00657856886344477,-0.00145573721035874,0.00587074223273953,0.00409457310342565,0.0112182862207668,0.00766776070524355,0.00542402843348522,-0.000725227892248381
"1469",0.0104705717535523,0.0115807678244608,0.00993350956308503,0.016281913171325,-0.00818739849908812,-0.00199575691469345,0.00109352156488107,0.0108001870839911,-0.00455550554989503,0.00181427353995822
"1470",-0.00889209836603599,-0.0122472018524079,-0.00765040520925264,-0.00526069768071835,-0.000735824554200626,0.000837049480058916,0.0067114625305269,-0.0111704353377207,-0.0208948085369804,-0.017022771955908
"1471",0.00204915583069609,-0.00377355036769988,0,0.0048077188192881,0.00564401072881293,0.00241636786788546,-0.00744181806876243,-0.000982337322203874,0.00387447710180266,0.00847457402154794
"1472",0.0078251670236511,0.0113637324119289,0.00220292894394114,0.00789490681541194,-0.00943504040508691,-0.00454259430976067,0.00218666807998491,0.00958669493005471,0.0188078605356334,0.0179027562684033
"1473",-0.0226638164709962,-0.0160514937927543,-0.0120879335929149,-0.0163783420811374,0.018146091605268,0.00838073123260052,-0.00498744183908795,-0.0126611252908436,0.00114252553561278,-0.0186646826118815
"1474",-0.0120241611529823,-0.010875385876179,-0.00444962061386045,-0.0125481648883712,0.0148391734519997,0.00443290765279336,-0.0101816322636803,-0.00838454405413003,0.00900954985255731,0.0014629624526632
"1475",0.000869198897281764,-0.00329873246686074,0,0.0019551603376371,0.00111241928908923,0.0000915310290610094,-0.00332334481806018,-0.00174074627506038,-0.00101195306232649,0.00803510311144295
"1476",0.000796373515276283,0.00193097827878441,-0.0100558207566921,0.00365862868250111,0.00166654904226315,0.000643898490579442,-0.0015877574480001,0.000248910543966252,-0.00220480267290191,-0.00471015522293972
"1477",-0.00347183960632891,-0.00330337353376975,0.00112875111443711,-0.00899161522824621,0.00332865539704663,0.00119395969275549,-0.00318083654393997,-0.00423424158257946,-0.00209012246205054,-0.00182014263204167
"1478",-0.013498582880925,-0.00938935133316776,-0.0124015031779604,-0.0154485906398831,0.000947782697934274,0.000275522516245408,-0.0194637747142488,-0.0120058291739553,0.000239335718515754,0.00291761361802267
"1479",-0.00169194256742811,-0.00111531427008815,0.0159820129086623,0.0034867378848018,-0.00197265533649771,-0.000458665646954293,-0.00439302108777995,0.00759493365860298,-0.00628217665598985,-0.00400002006035627
"1480",0.00493734398862555,-0.00558183299659643,0.0179776462464949,0.00297848169028536,-0.000869840466195093,0.000642263778981356,0.0114398370413165,-0.00175905235230367,-0.00126432057954895,0.00438110108307055
"1481",0.0202390969881938,0.0224529708755306,0.0143484095918061,0.0175698748745647,-0.00561832985946209,-0.00201784983219799,0.00937122173104776,0.0148503817821461,0.0119965634194428,0.0189023340870691
"1482",0.000431161364020216,0.00329383164439445,-0.0021762246516942,-0.00194553614549198,-0.0100276476521453,-0.00413584389076627,0.00624315455343116,-0.00247998590073761,-0.00285933171082775,-0.00677854216455243
"1483",0.0018679233319463,0.00355665906878988,0.00109068456989947,-0.00194912798043057,-0.000562205888389844,-0.00147613950033787,-0.000636712530511896,0.00124307576072891,0.00101558636128574,0.00431032299677248
"1484",0.0136250178395596,0.0239914417557368,0.0119823783531987,0.0163572086279857,-0.00096500779007469,-0.000554761835621642,0.00811868099694846,0.0144027660945421,0.0122344415401581,0.00357656282013474
"1485",-0.00212233285140428,-0.00213006535270888,0,0,0.00474978922188019,0.00166464481648387,0.00142130220672665,-0.00195824044157711,-0.00106130534130477,-0.0014254239409307
"1486",-0.00510470422958387,-0.00586967295338525,-0.00538198268502588,-0.00840731850671195,0.00392621009572025,0.00230803268507884,-0.00536125284471889,-0.00220758467685189,-0.00424946012952976,-0.00142760560061006
"1487",0.00805252455350325,0.00939338091955255,0.00108217847308434,0.00557172198130118,-0.00143645935717807,0.00128955556739707,-0.00174371240040705,0.00540816791731102,-0.0128030579715404,-0.00321664961115631
"1488",0.0046656044813782,0.00904003758986271,0.0118918237073187,0.00722715733181389,0.000159773858182,0.00101194228141344,0.00651105794674622,0.0083127553191602,0.00378258774333373,0.00681249553246777
"1489",0.000210862186729388,0.000790606582562026,-0.00320488360930238,-0.000478272694444559,-0.00271757855180443,-0.000184195118927755,0.00394453880616563,0.00193993811946136,-0.00675912218754549,0.000712314306763551
"1490",-0.00492388093352714,0.00368605173756364,-0.00428749926353489,-0.000478642300978049,0.000923940978135196,-0.000395346676670072,0.00282874728419502,0.000484108499620772,0.000481794631464139,0.00249106907856311
"1491",-0.00141392335525192,0.00524680581856107,0.00107656585590643,0.00287286292358679,0.00577550130424132,0.00174909433871062,-0.00125358086896088,0.00217685852142857,-0.0102931857493174,-0.00887467772603245
"1492",0.001769565039486,0.00182688257581409,0,0.0107421850317444,-0.000478670121833114,0.00082713350572261,-0.00266747353734031,-0.000482715521244237,-0.00182461381613697,-0.00107455759836994
"1493",0.00339221322435512,-0.000260782997411724,0.00537628546621538,0.00755807508062456,0.00215461823406016,0.000550829295068223,0.00881030309177677,-0.000241312706645846,0.00231540952703546,-0.00896381185338879
"1494",0.00302898861130729,-0.00286598318636921,0.00320855139450216,0.00304729909870494,-0.00923618297151207,-0.00284509016002921,0.00405497902040164,0.00942011302224488,0.00401218237082057,-0.00108533151390944
"1495",0.000421108965134698,0.001306551927994,-0.00319828951820844,0.00560887346468997,0.00442024244315053,0.000920747188879467,0,0.000239331960262046,0.00387502412509044,-0.00217317058423616
"1496",0.00680799429798173,0.00887267012537873,-0.00106920670276123,0.00511284958355507,-0.00760157255680438,-0.00193100026101223,0.00124248208121047,0.00311032196518202,-0.000904758729105781,-0.00181478263702284
"1497",0.000488671542153707,0.00439730313135134,0.00428233680047385,0.00300564689299843,-0.0116097557479509,-0.00423834793983802,-0.000620500697194326,-0.000715704749976953,0.000724479350117102,0.00472724539946046
"1498",-0.00613258348416956,-0.00283305513795251,-0.00426407658837935,-0.00437985488583226,0.000733848355910949,-0.00194256678551163,-0.00667477393005189,-0.00548929592618641,-0.0084454905363941,-0.00904819863907314
"1499",-0.00371549230945767,0.00490713267594711,0.00535325932910813,0.00439912240358509,0.00749914693592979,0.00222426940033627,-0.0012502804464759,0.00551959461441753,-0.00146005966599916,0.0062089023060381
"1500",0.011752081034724,0.00429222289462694,0.00958440859941656,0.00253564979558218,-0.0149673314803268,-0.00527219803302703,0.00625881678609774,0.00811453883596114,0.00188872838942511,-0.000725868225068038
"1501",0.0111288844221107,0.00875380880817045,0.0150336084790705,0.00698611584337216,-0.0101850266650363,-0.00390578678729636,0.0102626409321327,0.00639206428449524,-0.0143517390616426,0.00254264592044251
"1502",-0.00742924043979154,0.000765777852314908,0.0157565204699701,-0.000459266719449514,0.00331911728814549,0.00140048783672175,-0.00140233442201076,-0.00352833527760121,-0.00240621912134487,0.00362325082674775
"1503",0.00575195517944094,0.00586565731992406,0.0134434936708701,0.00597562937794849,0.000165918299551704,0.00065238674226431,0.0113906143364966,0.014400127630066,-0.0121219987368173,-0.00469318791637974
"1504",-0.00907710018715757,-0.00938105721731675,-0.00612254458206762,-0.0114233045810979,0.0109149538419155,0.00270218324073279,-0.00308554667749494,-0.00667187771372646,0.00375637647921812,-0.00181354069069395
"1505",-0.00308074669605585,-0.00204776047126831,0,-0.00208021258882496,-0.00179935595882319,-0.0010222735286326,0.00139254443521497,-0.000487252496968682,0.00180872573057145,-0.00327037887043391
"1506",-0.00421523855981742,0.00102591824609122,-0.00102678625943819,0.00301074426711812,0.00359666741441345,0.0020583114385011,-0.00494498342093197,-0.000973585633127771,0.000996164892173024,0.0102077748250822
"1507",-0.00134057232835783,0.00435567610913234,0.00102784163310399,0.00563566224019363,0.00335541542639617,0.00204470943218737,0.00124240457076485,0.00316852798159184,0.0023635091576284,0
"1508",-0.0108080732142044,-0.0142856914755879,-0.00718661934418729,0.00367454526270738,0.00570957479362133,0.00231895830778406,-0.00604959432646213,-0.00753202157044919,-0.00384717662330147,-0.00288700503424477
"1509",0.0169964736842563,0.0170807097329388,0.00827285949570933,0.0148742261335719,-0.017273796772671,-0.005274787079247,0.00920759477977406,0.0122400927658384,0.00921895517959803,0.00542888193349578
"1510",0.0256299179705479,0.0145039148175474,0.0246153130532256,0.0196168934855425,-0.0133684896631127,-0.0045586006914512,0.0162360322790014,0.0133011371721969,0.00709785194178858,0.00359966281133017
"1511",-0.00225910386417749,-0.0135440953261109,-0.00900881654300201,-0.00707675688843867,-0.0135496982788864,-0.00514037332696549,0,-0.0152746016769812,-0.0120733040641454,-0.00824960277536924
"1512",0.0043913684012078,0.00711918917394971,-0.0040405414994803,0.00200472435241905,0.0038998562535919,0.000469848737863598,0.006086427483593,-0.00169665754819492,-0.00471460926888234,-0.00433994176907604
"1513",-0.0027324005077356,-0.000757154821817263,-0.00912770626654535,-0.00755717985219717,0.000422669123452568,0.000563271110335606,0.00151240174733691,0.00315642962688556,-0.00629524424962291,0.00181617565745906
"1514",-0.00287727370135071,-0.00202137428893745,-0.0133060940934759,-0.00895868254896315,0.00658525070494198,0.00244016089771848,-0.00196291403539406,-0.00847075952674159,0.00708778178269132,0.00253807371799342
"1515",0.00254191486188016,0.00101267211899536,0.0134855338761326,0.00429381099322446,-0.000922749494106534,0.000561583660114495,0.00378250369988042,0.00488173153981597,-0.000435930498703718,-0.00144667207169502
"1516",0.00794923915844437,0.0174507900756165,0.00818838309982328,0.00877572496154255,-0.00277043091631834,-0.00290031874068652,0.00241171226992298,0.00777289516749557,0.00928401117564914,0.00362186399421871
"1517",-0.0000672775209601406,0.00422563002204646,0.00304550678002458,-0.00803016629054754,0.00892308687766485,0.00319032954033971,-0.000150270545544062,-0.00385647163402014,-0.00567970133793549,-0.004330618978589
"1518",-0.000680461018681244,-0.000742592003032949,0.00607296969320581,0.0042723583569011,-0.0027533260243533,-0.000374038134698496,0.00150406367399425,0.00435492407799631,0.00298022479796622,0.00652420086718264
"1519",0.000680924361165625,-0.00346783238967197,-0.00301826750774081,-0.00425418296276836,0.00460187900463649,0.00243267352503618,0.00465554049379624,-0.00192694535839955,0.00631425680450537,-0.00432122496650611
"1520",-0.000136234244481614,-0.00472273245937682,-0.0121088349302643,-0.000899562843790891,0.00208230532977982,0.00130684189671726,-0.00104649666651846,-0.000482942872436998,0.000553617132795337,0.00108497613651792
"1521",0.00646035471064121,0.0107389534694291,0.00408571415919545,0.00562700103852531,-0.00997350679273246,-0.00456796095207501,0.00224457846066728,-0.00217316931964118,0.00430379358021993,0.00433527532181133
"1522",0.00222983959069678,-0.00222374099229328,0.00406931518557041,0.00223786591463648,0.00772344041504125,0.00280972360478282,0.00597162080820302,0.000967729416909258,-0.00159173547872404,0.00647484275670118
"1523",0.00539329960431756,0.000247278417748742,-0.0101317195621293,-0.00156319367649349,0.00191578041480223,0.000840292530491338,0.00504634364195145,-0.00338462647242721,0.00355633094748486,0.00285914600816461
"1524",0.00160929653427733,0.00049540691187433,-0.0081883830998235,-0.00536775165805048,-0.00149670139313707,0.000466445576450925,0.000147639998018034,-0.00388173276504855,-0.00281047843600513,0.00106912297437733
"1525",0.000267689090018397,0.00569171622332143,0.0113518950970086,-0.00359801480028232,-0.00349744101393701,-0.00167830547778069,0.00118092646311596,0.00487085623299421,-0.0109675199021344,-0.000711914167553562
"1526",0.00562216359859824,0.0135335372770813,0.00714293087019024,-0.00338529127439413,-0.0137040535307879,-0.00663331169941517,0.00412931493137236,0.00581686869366149,-0.00477018962669051,-0.00213755737961818
"1527",-0.00119771379854783,-0.00194209655551891,-0.015197579343194,-0.00701985172689479,-0.00364362555287112,-0.00206886335692613,0.00102813111470446,-0.00578322841335566,-0.00224090266694921,-0.000357010471621177
"1528",0.00393088302450639,0.00510815863461445,0.01337454112965,0.0111744538031255,-0.0055272612469095,-0.00150780036239073,0.00190712054774589,0.00290824349671293,0.0043671597140813,0.00571428109331551
"1529",-0.00391549168471028,-0.00121019564210767,0.0101520654363589,-0.00473601123534928,-0.00170970114224955,0.000566357575088494,-0.00922513061974573,0.00338354432565202,0.00745386025672823,0.0113635906775538
"1530",-0.00246563677261691,-0.00411911548823396,0.00201023079447005,0.00203919976401834,0.00488250447508976,0.000848860450436639,-0.00576429375707577,0.00120403327872531,-0.00610398290765168,-0.000351118811761197
"1531",0.0102871743986703,0.0104623479157988,-0.00300907382538362,0.0065580555979099,-0.0129848858591542,-0.00339742310754176,0.00668961447777683,0.00384915473925784,0.00155086851521458,0.00386373583612265
"1532",-0.0112405197791928,-0.0276908848554497,0.00100590278740764,-0.0132554622744313,0.0128088896566203,0.00577652006064233,-0.00206736252223239,-0.0134196982671042,0.00340664608374075,-0.00349897458315218
"1533",0.0100973219696894,0.00693391660565768,-0.00301501104152291,0.00113865487922071,-0.00888730055039255,-0.00357755867304566,-0.00133208896436487,0.00607252870626862,-0.000246870370370411,0.00386237920578703
"1534",0.000728626447163538,-0.00270525568342606,0.0131048943980894,-0.00113735981891339,0.00819157685687633,0.00302323072603161,0.00177835308236141,0.0004826792500634,0.00265492702775694,-0.00139907150236718
"1535",-0.0013232868592522,-0.0120839150527655,0.00298512118005911,-0.00887954917336542,-0.0022236291010681,0.000470889798429575,-0.00473305000826096,-0.00627391048878301,-0.0033869265557418,-0.00385290912519543
"1536",0.00556467338678557,0.00848743244706318,-0.00396827891161644,0.00735120812372547,0.00385705553499527,0.000753747435478624,0.00995684771169025,0.0106846554249211,-0.00166824645744557,0.0038678114512305
"1537",-0.000197991489942373,-0.00594085753655715,0.0109560506889923,-0.000455981011356577,-0.000768966666314541,-0.00103490163059128,0.00102996410282552,-0.00336389486930688,-0.0115739921952223,-0.00350257911454177
"1538",0.00164731895021664,0.00821742169921524,-0.00689640444479245,0.00273777422747767,-0.00247775662445926,-0.0010365572382689,0.00587983516692892,0.00168758990981877,0.00118974329097821,0.00175744514794096
"1539",0.000854846737124104,0.00493940709049845,-0.00396827891161644,0.00500562847949992,-0.0081378553281769,-0.00348862549715123,-0.000438400374728976,0.00553565060641126,-0.00525358687381061,0.000350872390607826
"1540",0.000920653503454272,-0.00737311616119007,-0.00996016686119339,-0.000452677556651682,0.00906799355408139,0.00425756107299047,-0.00394759958392332,-0.00526550454054509,-0.00440111277457822,-0.00140306948977265
"1541",-0.00118225004641637,-0.00321841294767111,-0.00301826750774081,-0.00362390778320731,-0.00290994155263014,-0.000942019905847524,0.00117458411546356,-0.00433154598841612,-0.0163562418810391,-0.00421490567380778
"1542",0.00749449947225478,0.011177677044004,0.0151362399562276,0.00204571599275849,-0.00497821245681151,-0.00160296980905661,0.0068902782064324,0.0113580135682925,-0.00276061256935711,-0.00388012635360513
"1543",-0.0124630168994686,-0.0132649894585879,0.00298204376072975,-0.00884752896143393,0.00301937090810256,0.00217249139349129,-0.00844501493867944,-0.00740695278347714,-0.025043455545697,-0.0113313996413342
"1544",-0.0060792156706837,-0.0164301716558926,-0.0118927104598939,-0.0137331651097351,0.00584793634273195,0.00197895664419967,-0.00778259277632287,-0.00698114703246711,0.00779181843909371,-0.0114613456196369
"1545",0.00977289633275991,0.0151863647846833,0.0160480220933741,0.00440926662168128,0.000684190943848861,0.0012232351354724,0.00858397495606122,0.00509064990101682,0.00229331680950451,0
"1546",-0.0190268522342947,-0.0309152515073503,-0.0138203691086599,-0.0134008727423505,0.0196531155110411,0.00770396736023882,-0.0168747645655449,-0.015918955782969,0.00895597170062135,-0.00471015522293972
"1547",0.00684574868269894,0.00694639851315082,0.0190193637704128,0.00562064342987401,-0.00578170607049777,-0.00186477225695814,0.00880586079592471,0.0137253797618604,0.0121809320249042,-0.00182014263204167
"1548",0.0125977892506117,0.016607114810312,-0.000982488039925733,0.0109451854357145,-0.00295046065607174,-0.000467208688894272,0.00769339208808306,0.0108802642345929,-0.0105619894343746,-0.00619988201925725
"1549",-0.00197437927306987,-0.00276465169163975,0.00393316128781218,-0.0046072943769665,0.00185985448873227,0.00140187385277257,0.000146928059988838,-0.000717470829033839,-0.0101572551523531,-0.00440368522061918
"1550",0.00329752299062736,-0.00453621371646051,0.00979410816240267,0.00231462100042434,0.00544571329669785,0.00249427188557005,0.00190837399876953,0.00694090792532509,-0.00366011764705887,-0.0070032599178137
"1551",0.00532548291377188,0.00405043991411436,0.00581968402624078,-0.00946678965171266,-0.0052984202858597,-0.00232960519260139,0.00747265286366305,0.00499190448627851,-0.000918387550270405,-0.00371197812652269
"1552",0.00895835374149923,0.0115986719689709,0.00192870615363683,0.0121211477166445,-0.00287447935043805,-0.0010280491391369,0.00770802150542593,0.00402074318258072,0.000525292176126957,0.00931452061308158
"1553",0.00136159542689485,0,0.0125120826956542,0.00483657560658313,-0.00907329558696413,-0.00317885633452786,-0.00375252433783624,0.00235544532733067,0.00557810061759745,-0.00553713659489818
"1554",0.00181216242274362,0.00672960536613765,-0.00950570985025778,0.00275040495042345,-0.00770151097370542,-0.00384611014819292,-0.00362161373662095,0.00164535440497815,-0.00352407501204921,0.0066815377053342
"1555",0.00426433453239183,-0.000742411498885542,0.00479857444511067,0.00868584664554395,-0.0104347969150054,-0.00508570084964555,0.0005815153280464,-0.00351947835034894,0.000131017091741237,0.0029498120940703
"1556",0.00379552573274533,0.00322104737512485,0.005730216404771,-0.0054387225026955,0.000958667494635579,0.000473794164514318,0.00392330088522264,-0.00141291186092518,0.00183352751728982,0.000735284073664522
"1557",-0.00224315471689784,-0.0027167345208724,-0.0104460165635155,-0.0113921471906177,0.00722631596227963,0.00274349821773923,-0.00361839354907934,-0.00589467481066475,0.00784363004628963,0.00220426929571249
"1558",0.00141277750420565,-0.00247673528298287,0.00575803330775204,-0.0094490145653966,-0.00103737612603039,-0.000849371240636665,0.000290683372565992,-0.000474071401605269,-0.00343730457957969,-0.00513193244750831
"1559",0.00532396982443983,0.0139031185629406,0.00572517424143593,0.00418795937202909,-0.00302843998276248,0.000283306722655086,0.00537309166162325,0.0163736851062246,0.000130085900557519,0.00736920964057641
"1560",-0.0013203974544419,-0.00171412666837434,0.00948777930195432,-0.00903612344957649,0.0046865687958797,0.00349263986487158,0.000433465615631068,0.000281296923561047,0.00208229447277497,0.00219455661418477
"1561",-0.00551850950994126,-0.0139809607855373,-0.00469914698676854,-0.0112229719545273,0.00760190727328669,0.0032929053830788,-0.00274353672543415,-0.00726507768629692,0.0089610714285715,-0.00583944890513199
"1562",-0.0023229878269091,-0.00248770313983138,0.00566549490551549,-0.00709373452615458,0.0067729051369867,0.0030941358221992,-0.00709399684427248,-0.00613811445946255,0.00450506485696156,-0.0073420437609536
"1563",0.00698507173666907,0.00573583974795877,0.00751178511096762,0.00571545970786991,-0.01115546228834,-0.00383253505722192,0.0058324704543895,0.00356286777035209,-0.00454899404729647,0.00702653066856218
"1564",-0.00854262449199872,-0.0116540530493443,0,-0.0101822610077458,0.00964485106840529,0.00262790550399528,-0.00333429573207211,-0.00591693009772432,0.00566393144313371,-0.0044069196129316
"1565",0.00803324870571354,0.0102862899285232,0.0037277858553606,0.00382803662796194,0.000768007313723729,0.000373976113849261,0.00610903746312363,0.0128575263178659,-0.00447998080000001,0.00184431274578434
"1566",-0.0041775842562074,-0.015644742346657,-0.00928485269585322,-0.000953680034038618,-0.000938057514293433,0.000748905373223252,-0.000670458644384198,-0.00188091645468713,-0.00199291542283031,0.000736442796368086
"1567",0.00800255107223835,0.00479342948696604,0.00937186912011834,0.0143133627543379,0.00119533248337422,0.00102790714005874,0.00744059549252807,0.00894984624273509,-0.00334967781017526,0.00919792752690629
"1568",0,-0.0100428800275294,0.00464252955882816,0.00376271981180798,0.00852039846152075,0.00429585491449536,0.0015932363520057,0.00396832555960613,0.00413650462683246,0.00510390617331535
"1569",0.00307368112324502,0.00710125916234405,-0.00184838933703724,0.0021087807114557,-0.0050692961170733,-0.00185999327061914,0.00462693665626634,0,-0.00585738925169044,-0.00943056091566707
"1570",-0.00395740041945358,-0.00528828197206366,-0.038888596698521,-0.0107552581588561,0.00753165074481554,0.00265857425530558,0.00316645520469594,-0.0179028717222891,0.00142441569616869,0
"1571",0.00493450664035788,0.0108859223444255,0.012523839624667,0.000472909381782127,-0.00405432271825101,-0.00195396313256657,0.00258264582045831,0.0187023572203264,-0.0144824790131568,-0.00476013385914431
"1572",-0.0101388776216719,-0.00500868112998132,-0.00380571166638954,-0.011811899256527,0.00898925338467671,0.00419569859769453,-0.00529506999894735,-0.00720396555129454,-0.0111526410684805,-0.0169242426921778
"1573",0.00405824317006864,0,0.0410693643582303,-0.00286898143013248,0.0119361379014209,0.00399144315014888,0.0146739553222914,0.0203645750684263,-0.00291914689628192,-0.0011226621444842
"1574",-0.00449112602959045,-0.00604058049055201,0.00550467379214181,-0.00239763608417642,0.0201843126771701,0.00314364635213815,0.00269387348091166,0.0142237851629774,0.01676761672349,-0.000749411160418934
"1575",0.00676702930404405,0.000759455464496073,0.0100364844129619,0.00168239584720409,-0.0076532252037903,-0.00322577756569797,0.00933262475985264,0.00226188190341903,-0.00425360911267092,0.00299958406858414
"1576",0.00345704466192553,0.0055668319667328,-0.00812990741340436,0.0098369013342916,-0.00246139528746592,0.000370148125595771,0.000420646840766814,-0.00112851739679376,0.00775494196227822,0.00635520752959895
"1577",0.0122483511843356,0.0158531475802917,0.0209468515373987,0.00950334703969058,-0.0137360261479755,-0.00416024304532692,0.00588140641482471,0.00610027319022355,-0.0168905443299999,-0.00222887210996559
"1578",0.00327729332644888,0.00569699035098603,0.0115969140572698,0.000941481901095775,0.00191778247751695,0.00111393790560399,0.00487247594682372,0.0038180096580005,0.00199006965174142,-0.00409532978060922
"1579",-0.00244969496268221,-0.000985114550059452,0.0017635572251713,-0.0152834125743566,0.0148995856262744,0.00556339665449679,0.00581893390638299,0.0123041053635182,-0.0470043419992517,-0.0123363959983461
"1580",-0.0231739235664569,-0.0219428256535333,-0.00792239125649141,-0.0243553508447762,0.00869370776329181,0.00221291577133931,-0.0249312885519842,-0.022762282482362,-0.087808261642409,-0.0299015704037351
"1581",0.0147632256430208,0.0143687635848639,0.00976041426970631,0.0205582060529563,-0.00821207973377525,-0.00285196627723616,0.0158216754225853,0.0174128006390113,0.0113472319145111,0.0105344659073492
"1582",-0.0146119133959257,-0.0280817048644068,-0.00702982427539389,-0.0158273732201655,0.00664000714951296,0.00184517473545864,-0.0120987324789638,-0.0111135259435678,0.000527048180864798,-0.0146718133830123
"1583",-0.00625346135707683,-0.000766834707973896,-0.00707959256708202,0,0.00244331095409489,0.000552292622456374,0,0.000449586979022643,0.0107624599519254,0.0105799947329301
"1584",0.00869301432286074,0.00690881861798753,0.0106950563067425,0.0146199599950394,-0.00211186593247836,-0.000551987763686701,0.0115429300823835,0.0146031043859034,0.00871182407940818,-0.00232653110253789
"1585",0.00443840528915307,0.00482850549839142,-0.000881815371229888,0.00480291173418368,0.000732588492955655,0.000552292622456374,0.00139161375160368,-0.00221398494808533,0.0179374989448771,0.00310924862864859
"1586",0.0103088045474851,0.0171978859224107,0.00970865285166234,0.00478017754410343,-0.00349804593871295,-0.000643748738312966,0.00583663392211187,0.00199743818536735,-0.00739658480333205,-0.00619922233375714
"1587",0.000634114361900417,0.00795607420717848,0.00611892080499388,0.00594656579798336,0.00253080323060839,0.000460344078900388,0.0031776222439106,0.00442948546793098,0.0108853736526382,0.0109162716021534
"1588",0.00405352359575417,0.0051802235921774,0.00521313342637408,0.00898571401799031,-0.00431606141780128,-0.00110456814794424,-0.00123980097593945,0.00308705105389473,0.0235600933569451,0.0131122044342977
"1589",-0.00176608535249478,0.00294455428672968,-0.00259304880379163,-0.0100772628228746,0.00915984066043007,0.00359415621361858,-0.00455010086930197,-0.00395692676911275,-0.00508367559543632,-0.00570989639238018
"1590",0.00669811996161163,0.0149254820445135,0.00606565534603631,0.0104165421344098,-0.00364655232071787,-0.000367283479290381,0.0077570805685927,0.0134630630131622,0.00986444511065376,0.0133996281898012
"1591",0.00238560990977899,0.000482181490012223,0.00775203632564092,0.0142925183818192,0.000569140489955267,-0.000183819593064127,0.00975929974091727,0.00413730876685148,0.00330288819459823,-0.00755569810693069
"1592",-0.00876737396572536,-0.00578294564381832,-0.0111108735937188,-0.0108569376836294,0.010273118082897,0.0032661471478368,-0.0068062396788674,-0.00303635523813106,-0.011627113213501,-0.0178911993642445
"1593",0.00928744540393356,0.00484722654968994,0.00432125962797869,0.00794007478776471,-0.00129013583864845,0,0.00383740505790353,0.00478599152387926,0.00574018137807242,0.0127906433562244
"1594",0.010140655195477,0.0125421727457831,0.0137694278328364,0.00834087869349442,-0.0235772949071177,-0.00852834081973319,0.000819383604127477,0.00974240052625497,0.00119784387257416,0.0110984797220384
"1595",0.00254086449485125,-0.00214401690562793,-0.00424455638892696,0.00137893382452581,-0.00248060590392774,-0.00129418804110282,0.003956470744088,-0.00171529523406699,0.000422253513188808,0.00113548788016282
"1596",0.00506872965163097,0.00429701280147587,0.00170506451614361,0.00711316972837306,-0.00389638333473563,-0.00138969170968706,0.00584334784742602,-0.00536932796665979,-0.0124515587387221,-0.00340260002939397
"1597",0.00455106826903884,0.0125981290646164,0.00851057459203064,0.00774701058608529,0.00158148710835015,0.00120548132322695,0.00243172480357567,0.00539831328113283,0.0148169392072608,0.00455228966012333
"1598",-0.00281615847935313,-0.0103288083505114,-0.00759470445405763,-0.0072350752753555,-0.00257564068904559,-0.00018518976652826,-0.00512138453474653,-0.0124569903403183,-0.0115822611183781,-0.00037763835250948
"1599",0.00325360541617781,0.00403239387169751,0,-0.0077430545073407,-0.0107467180790081,-0.005651462238351,0.000270842340778232,-0.00282735293001179,-0.00859308299968875,-0.00453344997004712
"1600",0.000795475130133116,-0.00496093626553207,0.0127549453075584,-0.00918085502054711,-0.00766307559402513,-0.00176985325116752,0.00148981349501365,-0.00937858019167503,-0.00838118158820145,-0.00455409573522136
"1601",0.0103341519239739,0.00189956504031086,0.00671708744400479,0.00463290790795456,-0.0108618862950852,-0.00401384408146077,0.0052740122286361,-0.00440328147179292,-0.00447876205556108,-0.00343117818564065
"1602",0.00538607206222963,0.00402801732317348,0.00917437018870526,0.000230635101201582,0.00669127926055402,0.00262445184289528,0.00887785648362827,-0.0030959261248712,-0.0230751980708975,-0.00229530155362823
"1603",-0.004695003260203,-0.00330413992329148,-0.0148760807371786,-0.00345786652305935,0.0103974206358863,0.0047667107397158,-0.00319965977571179,-0.0015528810368558,-0.00401105979309735,-0.00115036996924256
"1604",0.00967695676510449,0.00710389208961182,0.0159395585119806,0.00439501432745959,-0.0126519287833768,-0.00539540662147064,0.00628651268782199,0.0135526394367327,-0.0225221052284915,0.0049904142640429
"1605",-0.0000599559923426529,0.00352726652571134,0.00660596921484147,0.00253355333439642,-0.00119596287514057,-0.000748626884063852,-0.000531412376003848,0.00548024445719331,0.0308994261364461,0.00649353610594772
"1606",0.00143780475321065,0.00234271858529711,0.00574256323812539,-0.0020677370795501,0.00786869733999085,0.00262141902714164,0.00465456888809723,-0.0089383664157292,-0.0165777833251103,-0.00569256107987448
"1607",-0.00741756048151532,-0.00864875471685123,-0.0106036337784639,-0.0110496599772396,-0.014850764200441,-0.00793567212074386,-0.024755220809306,-0.0217774876061739,-0.00707407408661687,-0.00458016862487476
"1608",-0.00289284301643655,-0.00495146190448448,-0.042044535421634,-0.00744863725632317,0.00473768390518781,0.00103520407952562,-0.0139811771517938,-0.0179899967036194,0.0202364632372829,0.00460124309412979
"1609",-0.000846266306112953,-0.000711120831067835,-0.0180721184362259,-0.00867759072561247,0.00137172622115012,0.000376374760540976,-0.00385445190417599,-0.0137388497235025,-0.00631458282211894,-0.00381682028174757
"1610",0.00598858540159597,0.00497964200557832,-0.00613512950310957,0.00544148965442459,-0.0253422492855889,-0.0117461980143644,-0.00995039849729373,0.00371425040195916,-0.00201846598454203,0.00919547400448573
"1611",-0.00649416980839324,-0.00542690974729476,-0.0167546880994722,-0.012705775531794,0.0112437814119848,0.00408853080842708,-0.0199607000484,-0.0168860955387242,0.0100381822594133,-0.00645409096761351
"1612",0.00369224305757654,0.00711760744966727,-0.00538124942925544,0,-0.00243206821381381,0.000094631775521048,-0.00954287997648673,-0.0115292456215491,0.013869279628135,0
"1613",-0.0143522020271276,-0.0209659723929581,-0.022542849003957,-0.0181125381442067,-0.00339610783875977,-0.00274500328144456,-0.0122232086889942,-0.0211855263566558,-0.0203364964228931,-0.0118455806241523
"1614",0.00550617393428099,0.00986520449778805,-0.0119925679918104,0.0148058512392708,0.00529856093738101,0.00144458268687964,0.00247494533846093,0.00437723829152747,0.0193398823079434,0.0123741931688792
"1615",-0.00480667580705574,-0.00381226957723713,0.0289449121700298,-0.0121983545614835,-0.00923487634705933,-0.00256315903418469,-0.0116178584356461,0.00750614471987054,-0.0093765954646764,0.0038197756843481
"1616",-0.0140011975188267,-0.0150680557417878,-0.0381125107867263,-0.0179176329316113,0.013805591044435,0.00485411981131079,-0.0107257253988788,-0.0206680799829501,0.00214455378672063,-0.00456618679793841
"1617",0.00905341034168661,0.00801355091707445,-0.000943271079539287,0.00838281431273891,-0.000606530283192686,0.00123135730031176,0.0187138683016803,0.00490825252905558,0.0074527373833313,0.00382265631848155
"1618",0.0127202746064268,0.00939525456786305,0.0387155622406703,-0.00513457418471241,-0.0178795243501401,-0.0077578503323088,-0.000583307124891186,0.0144076191733773,-0.0238042922713271,0.00228477333300514
"1619",0,-0.00167052808903945,0.0127272021740106,-0.0135166747598274,-0.00477193680193944,-0.00247900397157974,-0.00875274196813769,-0.0122773062618587,0.00495200333847534,-0.00379945755776012
"1620",-0.010315451648219,-0.0098018793047745,-0.019748630928825,-0.0189335526231873,0.0118983147867491,0.0024851647047528,-0.0153052319408443,-0.0216914738379457,-0.00515157525531462,-0.00877181068797406
"1621",-0.0082770302543913,-0.00120691858009259,0.00274749939992924,-0.00685633179777767,-0.0143031664860667,-0.00448120944349417,-0.0146465301893069,-0.00747371230518579,0.00750469043151969,0.00115427429577508
"1622",0.0152088035072824,0.0120859058649017,0.0237439057184301,0.0212219123506452,0.0156683965883704,0.00756615744795774,0.0304869771637544,0.0256019420721376,-0.00379884543761644,0.00653342551185299
"1623",-0.00627281718261152,-0.00740368527575408,-0.0312218812198769,-0.0157735589559027,-0.00236684233190232,0.00133095324003696,0.00250184919040852,0.00244750263714377,0.00515917432484025,0.00420005822399827
"1624",0.0077218180786478,0.00986520449778805,0.026703539229709,0.00915757108137183,-0.0052709830364932,-0.00237344098497094,0.00132129854793228,0.00366227308318079,-0.00490953681742734,0.00228141593051934
"1625",0.00790557649273138,0.00333571760402052,0.0170401911879823,0.00428572262057569,0.000529666074147395,-0.000570558776177066,0.00161322565712019,0.00997321036456045,-0.0122598411524305,0.00189678735838483
"1626",-0.0138169335336518,-0.0189979760031916,-0.0123456112433225,-0.0308734411931526,-0.0103281288455821,-0.0137105188750698,-0.0300101164492091,-0.0236030862430499,-0.0116552557460359,0.00151455709395831
"1627",-0.0247781357613819,-0.0326797496301096,-0.0410716398285941,-0.0448072328281519,-0.0164124916943522,-0.00453768508693797,-0.0390887902250323,-0.0434137462910712,-0.0535262900230122,-0.0325141227318189
"1628",0.00320999374789288,-0.00900907154090702,0.0363129066936978,0.0143709942386452,-0.0169589066858915,-0.0105694455630627,0.0117795186791905,0.00489224949821598,0.0117314322286639,-0.00625247726745759
"1629",-0.0126359921789592,-0.0154040286334264,-0.0278525573515637,-0.0203152346324078,0.00415135032244862,-0.00245053887223512,-0.00636436866275281,-0.019005352358738,-0.00895644120856198,-0.00432562145749138
"1630",0.00961423630855829,0.0118641450433667,0.0129390335611288,0.0212823164419464,-0.0089112068722359,-0.00117933794008229,0.0184346735242693,0.0177812598427312,-0.00371176470588241,0.000789878627295737
"1631",0.00990092650558849,0.00726355743720442,-0.00456194616802086,0.0157625207890999,0.00648875108144198,0.00403341849585326,0.0149571903655477,0.0104301413070758,-0.0420345181660766,-0.00276239324015415
"1632",0.00586983693558207,0.00463523708535574,0.0245787580794687,0.0200656674222264,0.0102228049081188,0.00538873637963855,0.0178489253252481,0.0198709348595683,-0.0197835392271182,-0.000395720742039196
"1633",-0.00409745501964776,-0.0066648439441952,0.00808614983939426,0.0057471354443428,0.00683728218291302,-0.0011696840528459,-0.00434656398074829,0.00961552789753872,0.0273417193834444,-0.00514652842086805
"1634",0.00586013803696162,0.0118708756515817,0.0124777078538023,0.00311707868244171,0.00201485442382965,0.000381176229920177,-0.00526850847802429,-0.00451131140796779,0.0169590796997812,0.00636692819458662
"1635",-0.000929473291423788,-0.0104564433424565,0.00704233465473769,-0.0178665818605667,-0.000633777896566823,0.000390625495655827,0.0116523741912389,0.0088117469388711,-0.00891599130477971,0.00395407799903147
"1636",0.000433915184222977,0.00128879696417683,0.000874235645459631,-0.00922736316653971,-0.0029906194085928,-0.00195254285353186,-0.00433818777628359,-0.00349401654095682,0.00574756337157267,0.00905876382185755
"1637",0.0107887005814729,0.00180169701962352,0.0131004129375549,-0.00638640697308734,-0.0340880448322384,-0.0168231967179581,-0.0105168017830461,0.00776346821467655,-0.0219480043390426,-0.00234196863799574
"1638",0.00570485226740547,0.0107913875215961,-0.00689636764254531,0.00133890384404833,0.00969335729280996,0.00586968869080362,0.00394774573162393,-0.00422440468558349,0.0120247781192235,0.00508608309389769
"1639",0.00719738430624939,0.00279613500057274,0.00520814531012448,0.0131050461310511,0.0010253004953289,0.00168092503869244,0.0127043906820092,0.00798601284984901,0.00928793390866134,0.0062280993616175
"1640",0.000363217225295198,0.00709748371972152,-0.00345430650098744,-0.00950356185586343,-0.00782142518177242,-0.00355419326878936,0,-0.00594200410240719,0.00273581488801655,0.00309481492883301
"1641",0.0136208235284865,0.0279388806029683,0.0294628173394231,0.0490404592729916,0.0117306273730649,0.0100080001524205,0.0276283206779262,0.0328763566100831,0.0272013318032576,0.00501346891729848
"1642",0.000417865465160983,-0.00759085164296125,-0.00168334029271122,-0.010670785508596,-0.000834543254314757,-0.000785278284194058,-0.0065394117855927,-0.00795748479614777,-0.000885391192617324,0.00383732509349644
"1643",0.00382078657730167,0.00444140859541808,0.00927470612024051,0.0102722758892468,0.00529129768496994,0.00314190312902163,0.00365663669897986,0.00607682260692521,0.000402827690393126,-0.00267588302880972
"1644",-0.0037469310913526,0.00122806480081739,-0.00835413462407975,0.00406716685150488,0.00341627666780897,0.000490064557443493,-0.00160321298319632,-0.00265763285201492,0.00571749879207606,0.00114992905154732
"1645",0.00256701808934467,0.00147204673455659,0.00926696323329801,0.00911411544478091,0.00184087064649829,0.00440178628841692,0.00525567824040052,-0.00314918040718337,-0.0125710546286417,-0.000765765091293669
"1646",0.00547749499940875,0.00857422935580243,0.00500825983278563,-0.0117915333187582,-0.0124928586674858,-0.00467512439726314,0.00624460316758357,0.00267326948426749,0.00559521569899446,0.00421458075059888
"1647",0.00177678795842851,0.0029147740549107,-0.00747507963978211,-0.0027923130298636,0.0158137054562308,0.00548002967828443,-0.00101046310110087,0.000969298760462589,0.00887024419207738,0.000763017835870849
"1648",0.00195070324802704,0.00484389615122538,0.00251054399534723,0.00992845592417546,0.00146529811567975,-0.0000974041597311404,0.00288917598860028,0.00508488609849023,0.0298137236846479,-0.000762436083540319
"1649",-0.00212362734698424,0.00168705522918611,-0.000834713821576627,0.0108393586651712,-0.00420663208909888,-0.00116749941228422,-0.000431864304010654,0.00048184902716164,0.00675264690321775,0.00152611420787818
"1650",-0.0036656172641002,0.00288750819650851,-0.00835413462407975,-0.0102242656853181,-0.0126717336391879,-0.00672414484971273,-0.0194552277477895,-0.0086684961184671,-0.0171922278903276,-0.00799996926074609
"1651",0.00243269788351053,0.00575804373938116,-0.0185342761272566,0.0057947986057485,-0.000372117397984817,0.00147127300790828,-0.00117594510796781,0.00364362736640333,0.0093347581737977,-0.00115205797759044
"1652",0.00106575304537238,-0.00238549227979767,-0.0231759545339051,-0.0022543614143179,0.00614071800451188,0.000881587512709281,0.00264884144944677,-0.000968367325002717,0.000854907917228864,-0.00615151468866593
"1653",-0.00307539256300438,-0.00382604624272109,-0.0219683520503358,-0.0125533745161952,-0.00730520923793399,-0.00205499140122445,-0.00792485715356184,-0.00823629179742569,-0.00240719057623229,-0.000386841912370151
"1654",0,-0.00336054411194509,0.00898461093266034,-0.00228817941574921,-0.000373038972691697,-0.000294241798009853,-0.00118373116378889,-0.0061066797076893,-0.00272441813089119,-0.0034830042132139
"1655",0.000712240752315463,0.00602143102746378,-0.000890460650768143,-0.00586139877329483,0.00363430958279598,0.000686755088858293,-0.0137735877813665,-0.00442348299779527,-0.00124879805060862,0.00699035586535879
"1656",0.0115581622487662,0.0100547645666818,0.0276294004909297,0.018200080418912,-0.0192683618876465,-0.00882615001671538,-0.00555646720491476,0.0118487357843153,-0.0105501563812922,0.00231393010372782
"1657",0.00169930455910805,0.00568875389511692,0.0156116315553585,-0.000251642604873759,0.0110101759637475,0.00851846361574782,-0.00437901775765093,0.00146388555955568,-0.00197456755410652,-0.00384769978730604
"1658",-0.00146245874369388,-0.00259270169804648,0.0025617140745906,-0.00629543792781184,-0.00769814550001446,-0.00314290961767816,-0.00060694447767462,0.000486906191689673,-0.00522320350408989,-0.00502117525665891
"1659",-0.00568249021733924,-0.00165396836227627,0.000851801383985773,-0.0126711986506385,0.00293299628394306,0.000295929278038454,-0.00349056000710979,-0.00146062368196598,-0.0137628961120818,-0.00815226196392715
"1660",-0.00324044736667084,0.00142044539343256,-0.0187233990044424,-0.010780370830044,0.00745209282183978,0.00364393157538401,-0.00411224648674025,-0.00658356911849656,0.00145197223963889,-0.00665361032499945
"1661",0.00366475813010236,0.0103992262106134,-0.00520379719143449,0.0192011272250223,0.00271499964975885,0.00147162648906218,0.00091762330921541,0.0112907821971069,0.0218284249403395,0.0051221547324638
"1662",-0.00288556906656046,0.00163710718691479,0.000871828350458959,0.0020363954578464,0.00158736361489353,0.000686282242729153,0.00947275855420338,-0.00169883731013665,0,0.00705608126312685
"1663",-0.00118128076239399,-0.00373647143275058,-0.000871068927872365,0.00940059558308892,-0.00680536519518515,-0.0019583391420529,-0.00817314856795792,-0.00705069567399352,0.0178937725217267,0.0120669074580908
"1664",0.00295652655067724,0.00609471032317899,0.00871828350458803,0.006040572233313,-0.0144563766398684,-0.00902663913704616,-0.0137339905178077,0.00171363976238936,-0.0107643998000311,-0.000384530976713426
"1665",-0.00512936585525914,0.000233217588825108,-0.00518573526885902,0.00325239323154891,0.00152403062269491,0.000890897972100513,-0.0021662658943552,-0.00097741995007905,0.00986380162617517,0.00807999927135161
"1666",-0.0139860454068882,-0.0051247301667271,-0.0139009451850375,-0.011471361044767,-0.0135042855871682,-0.00554007482169139,-0.0189175892211304,-0.00905333312837309,0.0208527286821705,0.0095419721382568
"1667",-0.00330569235609413,0.00210711640196637,0,-0.00857695749435483,-0.00347088339830415,-0.00387902827348807,-0.0230759466479586,-0.00074043398746082,0.00675829589553811,0.000378066669932675
"1668",-0.00639200233567072,-0.00887840207759238,-0.00264325967685353,-0.0188296871468735,-0.00870645560156313,-0.00429389810238867,-0.0135900194422538,-0.0113669084086631,-0.00429934372757068,-0.00113377136863213
"1669",0.00491592246926231,0.00353596343087847,-0.00883400487638997,-0.00181520731708229,0.00770962055630253,0.00541557203490672,0.023454342006191,0.00324949372773209,0.00333309610382138,-0.00189184165773648
"1670",-0.00616041094477171,-0.0112755804436938,-0.0142600684421138,-0.0233826622253877,-0.0109431971946916,-0.00628422601537526,-0.00208332145494339,-0.0174392675420095,-0.00286893173731062,-0.0011372096858524
"1671",0.00911534671354119,0.0125921977248018,0.00632903237831184,0.0162275796108744,0.0101830537386656,-0.000401405482456485,0.00562055748697232,0.000507138931050477,0.00560302082818853,0.000379579586898826
"1672",0.00337201229453288,0.00610042974417291,0.0170709596566356,0.0117801489108056,0.0108556494753291,0.00562347646577899,0.0116577402131697,0.00734955561907458,0.0157367369284953,0.00796658499444414
"1673",-0.00372075168332475,-0.00629665154143932,-0.0114840010155703,-0.0108665981739087,0.00498641634742492,0.00199713970477111,-0.00378840863547492,-0.00654085766036094,0.00407711656384513,0.00564542635091381
"1674",-0.0160842753435448,-0.0194789174906257,-0.0107238460716564,-0.02301866295041,0.0125939852495933,0.00568084143092973,-0.00301081970266548,-0.0157004341755488,0.00959765986558136,0.00973052179638567
"1675",0.00355091748906222,-0.00215436397626045,0.00271021710531438,0.00214174673761436,-0.00810288385837787,-0.00406303532747987,-0.00476794521151513,0.000771953915193802,-0.000292453382084168,0.00148263579272623
"1676",0.00158643113439472,-0.00263829147557737,-0.000901188243820683,0.00801518693605385,0.00797927004470966,0.000994777624159449,0.00159701738578732,-0.00128546495673598,-0.00614448070359619,-0.0103626668671772
"1677",-0.00316794057295644,-0.0108227670803879,-0.0198378618561539,0.00768583624855457,-0.00113098876346662,-0.00188856911588997,-0.00765292398568007,0.000514768211223426,-0.0091999708986521,-0.00299180861046588
"1678",0.00452244263163104,0.0143450293797505,0.0248391764768532,0.00631274278204219,-0.0141040579412488,-0.00567480670839327,-0.00835470724903054,0.0128635241596373,0.0133709929197368,0.00525124106240105
"1679",0.00827267600175308,0.00479385597242055,0.0152602273073033,0.0177729676250142,-0.00220667974765143,-0.00331065037267997,0.00712879904235031,0.00457207879307764,-0.0129012903225523,-0.00858201128343494
"1680",0.0012670300496469,0.000476875322934944,-0.00265251067899708,0.011813086161315,-0.013944362345208,-0.00764902469642192,-0.00852633817656645,-0.00177006667254687,-0.0182682825406718,-0.00225815504595728
"1681",0.000482002415553184,0.00643800790749616,0.00354617688207148,0.0147209256615468,0.00497340151794945,0.00608571280048809,0.018335170545158,0.00329290241880975,0.0147503558566646,0.00565820345158907
"1682",0.00957624814923097,0.0106607785461648,0.0256183648198507,0.0262630738404408,0.000485237765758928,0.00201574658167192,0.0197579406866581,0.021711885464589,-0.00178896765362513,-0.00637662282010609
"1683",0.00739676573357517,0.0128927753822412,0.00775193428949672,0.00755533972736067,-0.00698313070068901,-0.00462779716605655,-0.00125011688526133,0.0113663180119243,-0.0162049057962839,-0.00906001565387571
"1684",0.00313903334474497,0.00740549267210411,-0.00683751951668155,0.000725762885528836,0.00888854715650389,0.00505366228153226,0.00688376021034931,0.00464189990886799,-0.000303689073034463,0.00152390635694055
"1685",-0.0026565803255918,-0.00413509556470015,-0.00688475974170399,-0.011602529548285,-0.00135540961560021,0.000100801828257113,-0.00637042487681438,-0.00583651722377065,-0.0305998412437321,0.004944778001164
"1686",0.00224900765667368,0.00392180392689956,0.00519938417631205,0.00660298716115459,0.00387750599341152,0.00130690911001596,0.00218900119821175,0.00660467718674584,0.00117491973329531,-0.00302796768043412
"1687",0.00578757378468175,0.00597416143765428,0.0129310352024701,0.011175936633522,-0.00666348263359162,0.00220919278611187,0.00983004426598999,0.00801953521015064,-0.0107182209356907,-0.0125284973465647
"1688",0.0044627112622142,0.00137050318536391,-0.00425540572827832,-0.00216239116001926,0.00826363422644794,0.00200407287260274,-0.000772451210496627,0.00699130499367695,0.000395436940975102,-0.0103806785639978
"1689",0.0115740103807229,0.0253193894937807,0.0307693108134122,0.0418974376241923,0.012342380067413,0.012400052741663,0.0349464036372473,0.0277711649413752,0.0435572727272728,0.0217560449952168
"1690",-0.00167613104770947,-0.00489435140566452,-0.00497522106026338,-0.00531549188905167,-0.00590540687072327,-0.00345746756090681,-0.00388463379913007,0,-0.00196950996021172,-0.00380226857225308
"1691",-0.00699139612642619,-0.00558920215377201,-0.00833331930627246,-0.0223048100919977,0.00527000536898337,0.000991672653199771,-0.0172490535583808,-0.0112544103728105,-0.0287666110056927,-0.0091603372497493
"1692",-0.00462725040998935,-0.00382184803626051,0.00336141788891897,0.00356447828393947,0.00733884210297253,0.00376283352322826,-0.00641044280399006,0.000237212966185174,-0.00320409505473651,-0.00731889206234926
"1693",-0.00235408661393466,0,0.000837440663423061,-0.00852440668909249,0.0107864320899866,0.00364992354030091,-0.00660482605322099,-0.0018971874684065,0.000862414719033699,-0.000388042802127453
"1694",-0.00288999807418422,0.00225685053868618,-0.0025104513767078,-0.00764278614387581,0.00205907009379747,0.00275212108224676,0.0034336602941385,-0.00237504678187772,0.00885155071748245,0.00155269384311052
"1695",0.0038451285283061,0.000675611598614623,0.0159396723679954,0.00409150841296846,-0.00700606440316165,-0.00215668953286574,0.00606632418280317,0.00500004072614901,-0.00776451630057939,0.00775195220958547
"1696",-0.00459684681806505,-0.000675155455757914,-0.00743177905128478,-0.0117450184593179,0.00244590783321774,0.00137546194949922,-0.00371057673364783,0.000237120538909341,0.00923389929388918,-0.00499997149863052
"1697",-0.00532828426881171,-0.00653018304267816,-0.00831963616174847,-0.0113994986477234,-0.00150144259013518,0.0016675250264766,-0.0100868938254124,-0.00213175994233994,-0.00612551751472812,-0.00425197135461264
"1698",0.00791616977580589,0.00770617406369589,-0.00419446125447809,0.0198724506823325,-0.00303419701526175,-0.00222612071719797,0.0152061647920092,0.00688328825520768,-0.0280074675928559,-0.00659936835062425
"1699",-0.000944776657420765,-0.00134932626337358,-0.00505483436749365,0.00384876326547712,0.00151219130773628,0.00167042645546789,0.000617678480149486,-0.00117831798785673,0.0198250427747024,0.00976938764059976
"1700",-0.00922080170671802,-0.00495487170171172,-0.00762065615230845,-0.00383400707986847,-0.00160462946111772,0.00137418055082938,-0.0154322737522552,-0.00873297700088338,0.000944451455130668,-0.00154804612847681
"1701",0.00757675288116189,0,0.00170646268440877,0.0129898396957406,-0.00075616738743034,-0.00274433375977468,-0.00360502432108734,0.00309542003703256,-0.00511087435131308,0.00310081279751295
"1702",-0.00864468947197483,-0.00520597524735833,-0.0187391590709212,-0.00854869887457277,0.00406795397790871,0.000884480175840086,0.00440476813895363,-0.0113932551245587,0.00877262316266991,0.0069552021763386
"1703",-0.0116467291559202,-0.0102390412972611,-0.00347239310692171,-0.00958103200403826,0.000282515078115386,-0.000490722050858983,-0.0114331431390842,-0.00384111681307786,-0.00188026482200143,0.00345352149477884
"1704",0.000725134708132291,-0.00275862209656097,0.023519150284071,0.00749698216060835,-0.0080057672678564,-0.00176801961426298,-0.000316943672634462,0.00964056010470582,-0.0101255963873533,-0.00726575415014186
"1705",0.0215578754321537,0.0205164166441045,0.0144679932761642,0.0235238173180525,0.00161412242001524,-0.00216509502248585,0.0239303969244695,0.0181426535774594,-0.0145904685227938,0.0127119685621264
"1706",0.00644345276304903,0.00609894792735144,0.00167792377940001,0.00445584640259944,-0.000284770352045216,0.0014789789415075,0.00959624426181405,0.00281327520169783,-0.0134384730048719,-0.00532534128258155
"1707",0.0039936725498646,0.00291862061211412,0.00167513624140159,0.00583716276224044,-0.00805967758559623,-0.00334788352656457,-0.000306749500006864,0.0032732514103635,0.00187605223288823,-0.000382403970200285
"1708",-0.00725389769548901,-0.00268636818548884,-0.0083611190163132,-0.00974937818661881,-0.000669170281976994,0.000197691485484208,-0.00322044375965935,-0.00838940626757101,0.00732720821741917,-0.00344303107689314
"1709",0.0139659989817842,0.00718293555562655,0.00927470612024051,0.00796977352892436,0.0125309248141237,0.00484060081849091,0.0181537123232072,0.00846038386499415,-0.00153561784040357,0.00767759687630321
"1710",0.00668313273425514,0.0147093952544932,0.00835401904423039,0.00627930363834484,0.00906943289510775,0.0057019426069862,0.0154126161975292,0.0139832006867668,0.0314068072575133,-0.00533326056285455
"1711",0.00675456123390061,0.00636925546674316,0.000828604552449042,0.000924414822592423,0.0021534453573584,0.0000978258024066925,-0.00193448092443738,0.00873372059013144,-0.00447339514163236,0.005744925346165
"1712",0.0000571075054953685,0.0015277070154629,0.000827804007986988,-0.00161593882907751,-0.003176294526399,-0.000684758000320418,-0.00521847488428484,-0.0027345882544576,0.00102487191209888,-0.00228489091290041
"1713",0.0057914950855682,0.0126390519271182,0.00496287609754931,0.0097127667800867,0.0111525925545837,0.00694449485300996,0.0106416500462583,0.00525496174780238,0.0185855484662416,-0.00114502251469084
"1714",-0.00478879856109771,-0.00602550684524195,-0.0205762090047192,-0.0233622006975779,0.00389297130334509,0.00174843587556328,0.00207612175382654,-0.00659071716835458,-0.00502546791481284,-0.0152846645628761
"1715",0.00332238901312976,0.0073609259099976,0.0100842071628604,-0.00211074526170762,-0.00387787484784452,-0.0020360156328536,-0.000739849049478991,0.00205870837636346,0.00940237766100904,0.000388042802127453
"1716",0.00456747418073933,-0.000859772519551827,-0.014975032021709,0.00470036708814048,0.00370781409568899,0.00174928686244913,0.00977480990353441,-0.000228257711755275,0.00431110874416207,0.00310321811263736
"1717",0.00159126233986617,-0.00408691783636539,0.00337828789945305,0.00584776208281812,-0.00341721104153159,-0.000969731542251662,-0.00689374846398394,-0.00411040591222966,0.000766449445307904,0.00386688312838346
"1718",0.00533419744304386,0.000648058630437598,0.0075757533410139,0.00325609025050366,0.00129771930569023,0.00135857839953335,-0.00841820368466362,0.0011464208153007,-0.00605081197994506,-0.00269645895743109
"1719",-0.00496695341068454,-0.00366934131024177,0,-0.00556330971407748,-0.00601521613068068,-0.00261769548859547,-0.00729791744870789,-0.0084745030925113,-0.0013099945654621,0.00308999375752017
"1720",-0.00283655496955459,-0.00498256539859021,-0.00501262871665498,-0.0102564520467331,0.00214150329710705,-0.0011664675616494,-0.00720187854653753,-0.00323399686344583,-0.0143519129158065,-0.00847131645656707
"1721",0.0023894202433159,-0.00631396941287843,-0.0109151045590405,0.000471024852145119,-0.0108248725466759,-0.00554628316462735,0.00634706068114732,-0.00324445717262822,-0.00618444506316651,-0.0124271349969011
"1722",0.00351862295737471,0.00591587228183776,0.000849002971733404,0.00612073896584109,0.00094195811858655,0.00196021100171184,0.00135172587658694,0.00278998754897675,-0.00110278852546963,-0.00432562145749138
"1723",-0.00316708923672326,-0.00936627465644813,-0.0084818655471447,-0.0201217802099829,-0.0119481857557827,-0.00450055394042093,-0.0151470784473773,-0.00765139441805429,-0.00197145338650662,-0.00276465649222335
"1724",0.00510600464940314,0.00945483120231949,0.0136868306564424,0.00310395230403859,0.000476276293902123,0.00304648952817921,-0.000151904680967041,0,0.00505688219116451,0.000792149946476695
"1725",-0.0126436498257974,-0.015465070467779,-0.0185654906184489,-0.0180906468869231,0.00847031994385716,0.00264573257820899,-0.0121843908119185,-0.0135511717907881,-0.0081760457903155,-0.00712309554301804
"1726",0.0134912233320315,0.00553097805901825,0.00773879441853786,-0.00218209430706484,-0.0240655122219087,-0.0112370500810279,-0.0134131829790171,0.00450025348486705,-0.0149017512713459,0.00557991813609582
"1727",0.000169304974336537,0.00308031374899875,-0.00170658072969698,-0.00510185632187232,-0.00377172109217438,-0.000494089174967294,-0.000781477602735836,-0.000235804709581733,-0.00329897009413405,0.00435987023310913
"1728",-0.00202995697651231,-0.00592257090591186,0.0128205146396987,-0.00537255357740329,0.00465941390705349,-0.000889963708591845,-0.00344079944324727,-0.00165072589621562,-0.0114636793865259,-0.00670879114630474
"1729",0.00802417162164337,0.0044132948327138,0.00759500315307493,0.00171883709425935,0.00367162646223451,0.00415651211415335,0.00706222942080359,0.00118095467556589,0.00326664769130214,0.00437042702655299
"1730",0.00498966939554535,0.0024165190128973,0.00837512502979609,0.0161763221232361,0.00616083474117235,0.00482866302410501,0.00794758299302001,0.00802280510050624,0.0115588036069809,0.0043511245202319
"1731",0.00435062096317518,0.00416383917135721,0.0141195821076014,0.0190546557783398,0.00200909891233181,-0.000784041568771099,0.00247361364834697,0.0124060103928125,0.000402373873075623,-0.00157540193747197
"1732",-0.00349898689398742,0.00240080209590987,-0.00163807142312289,0.00899392584692538,0.00601507674423352,0.00353306288436239,-0.00694008615319675,-0.0034681163135869,-0.0114221203346203,-0.00670606351599057
"1733",-0.00217378256374046,-0.00239505204992851,-0.00574224828486836,-0.00609898552417576,-0.00759281773863185,-0.00371651620564217,-0.0076099527362985,-0.00719220730170389,0.000406794134958588,-0.00158862234773016
"1734",-0.00312797574269519,-0.0104758061977032,0,-0.0136888444427538,-0.017023716960212,-0.00549781516041792,-0.00876358591289939,-0.0100496199331559,-0.0230174385445491,0.000795534102772777
"1735",0.00806875580758382,0.00992514195437089,0.00412549658987782,-0.000957125435392392,0.001654396177168,0.000888647580564506,0.00536781175888645,-0.0016521533124173,-0.00149850978608446,0.012718632235597
"1736",0.00500250303088379,0.00502293061648729,-0.000821773019853089,0.0071853871050096,0.009324636070285,0.00286032762923893,-0.00298342505703675,0.00118217094448081,-0.000166783388914737,0.00313971495238485
"1737",-0.000995384126099674,-0.00173867933385607,-0.00740149386062294,-0.0128416456783353,0.00288710897558042,0.000785943925406984,-0.00425271876474997,-0.00661308569464159,0.00450301041532697,-0.00117365263192004
"1738",0.000276543896056358,0.00152382121820271,-0.00414222040619749,0.00337263281551858,0.00374257574356962,0.00216220368903364,-0.00284734101158668,-0.000713068494845093,-0.00531295870258142,-0.000391771302957644
"1739",0.00243517860892917,0.0036949663322956,0.00415944976388816,0.00648238938648338,-0.00172104743494128,-0.00225510661994788,0.0103108247968431,0.00499630370999071,-0.00300451510599231,0
"1740",-0.000662418373734375,0.00346471371518486,-0.00082830653448851,0.0102575713250397,0.000287606233707383,-0.000589748567991988,-0.00926367190859001,0.000473375237840523,0.0103800268741003,-0.000391844188296631
"1741",-0.00259652660639664,-0.00798428756757363,-0.00248757611493755,-0.0210151345879274,-0.00777836802224463,-0.00429467036265774,-0.00522973698409102,-0.0134879167840597,-0.0258491721420673,-0.00117599337105756
"1742",-0.00432082696809077,-0.0100066291041776,-0.0041562686348624,-0.00337670046623118,0.00367732462844028,0.00178083466337275,-0.00111513604005553,-0.00407797863070336,0.00323181658051008,0.00588701097795474
"1743",-0.000111004325971775,-0.00549340805262788,-0.00751260916758756,-0.00121024589224372,-0.00954535050922545,-0.00454259537094559,0.00223290295962553,-0.00192650506758107,0.0169549001098246,0.00195089246041613
"1744",-0.00439575958316485,-0.00397693100750562,-0.00841022858947127,-0.0058152799830804,-0.00282326143544809,-0.00247947404912308,0.00111395405377812,-0.00506754047488789,-0.0138379127529001,-0.00116836855358804
"1745",0.0111769216273787,0.0135314278478669,0.0127225284285621,0.0221788872351829,0.00478368317510691,0.000894598090539267,0.00778892145753152,0.00654873959250346,0.00211327129044969,0.00350880445250534
"1746",0.00254224131950931,-0.000437737140972727,0,0.00143067734821378,0.00233183260218084,0.00119261169429952,0.00646686630721161,-0.000963834115017104,0.00986923635927694,-0.00349653579214948
"1747",-0.00358303554419093,-0.00394112322734064,0.00167513624140159,0.00047618367382829,0.00717351914994047,0.00416802936663085,0,-0.0024121120416799,0.0175409203346064,0.00311894620786823
"1748",-0.0112309662055105,-0.00681480751162811,-0.00919748309266799,-0.022132386347068,-0.00770001004252918,-0.00385452782964701,-0.0216267132702344,-0.0159576362610973,-0.0078804711869972,0
"1749",-0.00330135737808201,-0.0108456199937736,0.00337550766235628,-0.00584075419881425,-0.00378224896940171,-0.00287688600417635,-0.00672751746140698,-0.00491406939907235,-0.0212642725362876,-0.00932762588406888
"1750",-0.000112109101982005,-0.000447532130515294,-0.00841022858947127,0.00244805840814188,0.0048680718120071,0.00149239908710075,0.00403154153573704,0.00197550707721383,0.0092146080884723,-0.00392313431467806
"1751",0.00623186656309271,0.0123126438929264,-0.00593732231121935,0.00659339637593104,-0.00368201906469412,-0.000496586454150849,0.00112441260642426,0.000246438614487809,0.00259679182267036,0.00315080387494393
"1752",-0.00318042367117954,-0.00457720944830442,0.000853042469743492,-0.00873391890871733,0.00447361461474949,0.00318014831375346,0.00529436223512247,-0.00812998900622053,-0.00868911339812661,-0.00471136123717364
"1753",0.0170726396270175,0.0156250678515926,0.0195843596584198,0.0199042973570234,-0.00503460568673464,-0.00376475790084452,0.017555032759945,0.0116741212466316,-0.00876528430231294,0.00197235968110299
"1754",-0.00115570429324852,0.00307697820290587,-0.00842440523321475,-0.0184020221298921,-0.000973201437136417,-0.00417671116639817,-0.0122334003848724,-0.000491130578065491,-0.0237224808798361,0.0023622536040393
"1755",0.00581641500306818,0.00328649997859531,0.00339834018932472,-0.00147985747201518,0.0153889516617733,0.00309574198218776,0.00778026471258819,0.00326213871422731,0.00975441560703727,0.00785547348507354
"1756",0.00534300345481298,0.010919357534348,0.00931406896759879,0.00741104440324669,-0.00565921884500031,-0.0031859480152705,0.00141550526549317,0.00825426439615118,-0.0031913230431031,0
"1757",0.00219122743358402,0.00691319724930439,-0.0134228359550707,0.00588526475980555,-0.00800686315815546,-0.00389511272645382,0.00174683969065126,-0.00173662697034993,0.00458594791035738,0.00311765026524369
"1758",0.00508414021573378,0.00493435835365585,0.016156482065093,-0.00853253166551993,-0.00385389632031807,-0.00086379700696626,0.0011097355163423,0.00372776395948216,0.00551248932838044,0.00155406033549488
"1759",-0.0000545283680146724,0.00533736705027787,0.00502103894533423,0.0154905634686311,-0.00284015541934879,-0.00060314976292275,0.0012665914581742,0,0.00325513968228774,0.00271524598323292
"1760",-0.000163037145188172,0.00339772294065455,0.00915905475772538,0.00435820754362815,0.00687565412849334,0.00271564726934415,0.00079075683705665,0.00940836781253185,-0.0147712086380325,-0.00580270831542484
"1761",0.00473264905078929,0.00423289818828421,0.00164997712953463,0.00771484612167206,-0.00634110493312812,-0.00451376041987439,-0.00316035012341331,0.0105466963598175,0.00632640615587476,-0.00155639897877735
"1762",-0.00958356316129172,-0.0229716857382819,-0.0164743563555104,-0.0385167687538027,0.00304314231422054,0.00392944780235549,-0.0015854328284004,-0.0189320883082098,0.0161901218690117,-0.0144193330254777
"1763",-0.000164148993750945,0.000862960684752112,0.00586270400886524,-0.00174172042647325,0,-0.000602332539816564,0.00587491175072175,0.00544289578639012,0.0109322118644068,-0.00632664688813733
"1764",-0.00289786410838289,0.00172422747178036,-0.00333068177587947,-0.00947162789594769,0.00420883959447149,0.00281236379833372,0.00410417782644656,-0.0034451185756581,0.00176040739575489,0.00119377599891823
"1765",0.00614197097529123,0.00709963104823497,0.00417735713167433,0.00427763815860294,0.00253393293599768,0.00160203617285415,0.00345845017308788,0.00172878421499378,-0.0056903765690377,-0.000794901731337117
"1766",0.00021772512994267,-0.00170909997124435,0.00166386382097339,-0.0032570721602414,-0.00272183553689509,-0.00489914565176375,-0.001566529910352,-0.00419030132025022,-0.00589123884867859,-0.00954649111203931
"1767",0.000653971183518731,0.000856025767816071,-0.00332238242692806,-0.00527915881610541,0.00584906974896482,0.00261249291216981,-0.000470786676267765,0.00173262291237841,0.00287839477958696,-0.00803205995609246
"1768",0.00272281115505169,0.00962159382112371,0.00666675469838185,0.0176900769625659,0.0119209316087625,0.00841872138655053,0.0119309492341502,0.00716572903156787,0.015195027985776,0.00647764372042814
"1769",-0.0133048423079348,-0.0084711242005906,-0.00662260342587684,-0.011919513575515,0.00498019045146325,0.00288200610242351,-0.0065157112018388,-0.00662408375018064,0.00631959909663071,-0.000402247119002164
"1770",0.0108975682261625,0.0128149909229103,-0.00250009308552912,0.010806914832306,-0.00457439592135578,-0.00376622659220338,0.00624625546574475,0.00419851331431453,-0.00933728332516814,0
"1771",0.00538985889281807,0.00421774917933382,0.0075189170527592,-0.000248676275743098,-0.00105309287740618,-0.000894674663151296,0.00465545121731714,0.000245766759176869,-0.00191838353422624,0.00281690432515114
"1772",-0.0012995874004057,-0.000209956610136786,-0.00331662251152542,-0.00547121515160165,0.0067089255764925,0.00278748514661253,0.00231682321052595,-0.0012290359800704,0.00108638639189751,-0.00160515579427789
"1773",-0.00422956700128185,-0.00483101887592197,0.00249568149589741,-0.00500144410994274,0.0041887215914731,0.0023829870253278,-0.00323609370461708,0.00221545815062152,0.00951664571736677,0.00120581268813291
"1774",0.00294053042570286,0.00548753134695801,0.00165972168427775,-0.00150775113746604,0.000758588391402304,-0.00108927589143226,0.00695712994452125,0.00343912755640563,-0.0101711982138428,0.00240863827526017
"1775",0.000652006386310244,0.00125941132504148,0.00248561662625102,0.0133400330561615,-0.00246304490935634,-0.00277658905738409,0.00261049093422372,0.00416114442764393,-0.00426060996476041,0.00480578379051
"1776",-0.0081933803890436,-0.00167703621381354,-0.0198348121820553,-0.0245903452859302,0.0141499761106016,0.00676125901443192,-0.000459620862911514,-0.0107261338332463,0.0218139018069652,-0.00079720148395801
"1777",-0.0213363032958803,-0.0317092879170057,-0.0151770523348445,-0.0262283736580906,0.00646135292086591,0.00404886247004388,-0.0147081682991647,-0.0197140777501844,0.00410542734128061,0.000398959814302602
"1778",-0.00491902574265513,-0.00542202168270289,-0.0128424502933567,-0.00392274582579388,-0.00697822614169796,-0.00304856010883958,-0.00606421244286059,-0.00351932275731481,-0.01087580332917,-0.00677829885603132
"1779",0.00595490911733032,0.010902874259501,0.00867311158203132,0.00630089483621843,0.00243620919865961,0.00147980195958741,0.0101686335918805,0.00983826026191981,-0.0000826884927470628,0.00481735918529047
"1780",-0.0096054547269504,-0.0138048994695855,-0.000859900778935718,-0.0143490338441313,0.00822475608931095,0.00472883652116485,-0.00464592459848567,-0.0102423300495893,0.0125672099024525,-0.000799030209567286
"1781",0.0106004926372127,0.00393679481998976,0.00172097445265562,0.00926427781398931,-0.00287359371812734,-0.000980289235322895,0.0121364792061904,0.0070673824676506,-0.0220462478807361,-0.00399842815131779
"1782",-0.00585833784827938,-0.0137254264130815,-0.0266321894469745,0.00157339101224196,0.00669389860081071,0.00392605762779574,0.00307427973584695,-0.0105264207220075,0.00267177931047291,-0.00120436045501515
"1783",-0.0225051595945247,-0.0203225140704832,-0.020300166346488,-0.0282796919684274,0.0121848748844156,0.00543566951744134,-0.0145592193004671,-0.0167173254910392,0.0102423519108119,0
"1784",0.00700444647111387,0.00901909764458209,0.000901132483273948,0.0202103240044194,-0.010611245180131,-0.00301996778968983,0.0104198746612645,0.0118497820628358,-0.00272009561490272,0.00763659306640951
"1785",-0.0012541507810091,0.00402244963123244,0.00180004910573128,-0.00369794103753229,-0.00924552861865469,-0.00361485633276293,-0.000308066641493743,-0.00152745031358559,0.00247956860037313,0.00199447064194791
"1786",0.0131870236848584,0.0213667269439997,0.0116802334956105,0.0209436636374025,-0.00429271222978633,-0.0018632018231366,0.00739046268540244,0.0137678040827149,-0.00041225986963267,0.00398087837775551
"1787",0.012395841121956,0.012421079702134,0.0159858724133979,0.00571297687765493,0.000843761285098221,0.00265261005512452,0.00672480625196936,0.0125760216481368,0.00767073585732003,0.0114988169728101
"1788",0.00183654503715558,-0.00258310370370662,-0.00437079147033703,-0.0111025689398977,0.0028089176091286,0.000489634849117015,0.00910895870784256,-0.0057131413080137,0.00613898675843472,-0.00548796906493509
"1789",0.0109438690827774,0.015105909111057,0.014047402853854,0.0216711016917601,-0.00578908365636754,-0.00440648916029773,0.00345990867401746,0.0174871997763633,0.0117149611408225,0.00512409213369813
"1790",0.00049479278079323,0.00276359674195947,-0.00173157114081068,0.000255515701197195,-0.00516627865873398,-0.00236104893495559,0.00060009643877601,-0.00147350893758391,0.00056287390991594,0.00196075756439518
"1791",0.00516255623420525,0.00678394572701713,-0.00867301630975614,0.00102191857587663,0.00566472983388611,0.00473302880951776,0.00389533373690831,-0.000491278314374233,0.00851882986418051,0.00547949829681849
"1792",0.0055189592932734,0.00547461871072863,-0.00437444781209861,0.0122512335066107,0.00056329747363093,-0.000687246466676616,0.0040300243680802,0.0036896599609757,0.0132281777548517,0.00350334094595328
"1793",0.00119533457877141,0.00607356540452497,0.021968434938447,-0.00932949930542448,0.00225205273089468,0.00245526501735638,0.00594613343731032,0.00955864799571127,0.00196618164425977,0.0143521342519306
"1794",-0.00662160004056744,-0.00666126285837132,-0.012037973346854,-0.00687193694439225,-0.00421289777822687,-0.00195928188894012,-0.00029542352120937,-0.0024274385774451,-0.00886974083406999,0.00267682779140133
"1795",0.00590089021151297,0.00586756618006889,-0.00609221837615492,0.00358800816403715,-0.00244400299401393,-0.00107954014424894,-0.00177399002256895,0.00803098443809236,0.0105329930434701,0.00190703312623652
"1796",-0.0011407307585003,0.00166685290582569,0.0078807713886615,0.00689463201147733,0.0052775797272131,0.00127736915171983,0.00162895785027306,-0.00193114732643462,-0.000156708466406141,-0.00266463921158044
"1797",0.00554697009199367,0.00665542287086551,0.0112945193056191,0,-0.00253140440513766,-0.00098149301401762,0.00162643819380337,0.00241882801603155,0.0110519123522197,0.00419845517025497
"1798",-0.000378697538206851,-0.000826390644169006,-0.00343629509873367,-0.0114124369315098,0.00892871502885217,0.00343811323637011,0.000442648879620755,-0.00241299140481899,0.00170557400939697,-0.00456098027062002
"1799",0.0000540505803139357,-0.0047560958093017,-0.00431033972535777,0.000769643570279976,0.00530996041745291,0.0029367103281932,0.00280302118598419,-0.00362890328543086,-0.00851331894131058,-0.00267273931650935
"1800",0.00524782075030594,0.00540201989152056,0,0.0189692573666882,0.00546648696459173,0.00117133916126799,-0.00102975020528717,0.00194266098861773,0.000702490042131743,-0.00306282394495516
"1801",0.00252900110250764,0.00289321179485857,0.00519473719925823,-0.00679252792586793,0.000553203491120424,-0.000975169954046784,0.00662727855097667,0.00508819430819596,-0.00452413427123555,0.00345609488391885
"1802",-0.00703208478671002,-0.024727177680151,-0.0232556412246436,-0.0177302915576182,0.00667538467105611,0.00494634630495061,0.000731742173019523,-0.0106072481077197,0.0209214068111252,0.013777356550581
"1803",0.0140557388877309,0.020283371371127,0.0255731977922884,0.0170188944125849,-0.0150416905616789,-0.00768428062613569,0.0122806344335695,0.016081935033075,-0.0123570503223529,-0.00377495795619198
"1804",0.000906325609104863,0.0012422612932097,-0.0111780017281133,0.000760899137216553,0.0021415336921129,0.0010787507462211,-0.00129978607932235,-0.0031176115124476,0.00163200195387003,-0.00833649397690217
"1805",0.00229004513861897,0.00868671854690772,0.0191303814570809,0.0141880258238427,-0.00984959434931176,-0.00430867803198431,-0.00477224185117076,0.00793812010706563,0.00993094118962645,0.00917079873772564
"1806",0.000425220216266009,-0.00676636732518721,-0.00682612226336032,-0.0127404587740887,-0.00628726194572893,-0.00432682499338544,-0.0113338632009318,-0.00119331563177261,-0.00829685808245906,-0.00454367128187516
"1807",-0.000531182815156961,-0.00639965808699117,-0.00429552812608569,-0.00683214464554072,0.0014165200827696,0.00108644306985273,-0.00367433106738735,-0.00931859702531901,0.000309931065455959,-0.00836828159099012
"1808",-0.00494263817544527,-0.00498645700951406,-0.0103538086391934,-0.0112098644499865,0.00264075323146007,0.000986567287405871,0.00545793104005998,-0.00651283586208995,0.00565318649217117,0.000383577422433889
"1809",0.000267277844528291,-0.00292351817172676,-0.00959006777714189,0.00206103867050556,0.006959958398427,0.00394265706538088,0.00220077633713878,-0.00534078298233887,0.0146310949127437,-0.00268401243046767
"1810",-0.0112134123820762,-0.02157048165579,-0.0167251778264309,-0.0179993921395001,0.0134503851114542,0.00589002552655638,-0.00322056818880601,-0.0126921123212573,0.0034153917507358,-0.00461366569400934
"1811",-0.00280807641683223,0.000856030068780989,-0.0116385028428202,0.00549871172457905,0.00018419304099937,0.0000977250098852522,0.000293601224904627,0.000741432020090915,0.00673170677617474,0.00540753876743816
"1812",0.00904358733840627,0.0130453541950233,0.01086969689379,0.0122396249363321,-0.007463709426204,-0.0040014239480054,0.00161508621774842,0.00914052473755422,-0.0109692481907178,-0.0111410364454776
"1813",0.00713818697079316,0.00865526450420884,-0.000896090643081271,0.0138922608468424,0.00362057060506471,0.00244981138907208,0.0043973510507278,0.00538546706180298,-0.00774843518496227,0.00505051615747321
"1814",-0.00532905034850362,-0.0146504454250187,-0.00538126753103341,-0.0213140827423643,-0.0077706975199513,-0.00928543948696603,-0.0176590609235729,-0.0112005304635125,-0.019369155541615,-0.000386463282109228
"1815",0.00583971728028421,0.00127439146476638,-0.0144272567611762,0.00440748655482404,-0.00177140875724935,0.000197482245725356,0.00133712984215628,-0.0123121184132521,-0.00179557348100801,-0.00464046671164819
"1816",-0.00387868170735994,-0.00318194896424873,-0.00457483579759332,0.00619520481059088,0.0108341076854326,0.00187382352425569,0.00816020224541458,0.0017062341816807,0.0047708430723381,0.000777070152832904
"1817",-0.00413537772653361,0.000212873110862155,0.00367663335574586,0.00974860343881101,0.00711456414248279,0.000394147944685397,-0.00588627946142206,0.00325670036026393,-0.0178251808373535,-0.000388273345873769
"1818",0.00474560066415375,0.0129786616317988,0.00457882452032443,0.0114329634531083,-0.00376156169298103,-0.00059049050744997,0.00732229184977751,0.00998761356338718,0.0018228245363765,0.00660197167429399
"1819",-0.00719235006364405,-0.0018903071352383,0.00729271209442195,0.00226084906970514,0.00782770740773975,0.00423418826579014,-0.0111492938047263,-0.00494459165353811,-0.00791076630295806,-0.000771634106060737
"1820",-0.00210800249640775,0.00273568176848604,0.0144794790417586,0.0130324085868923,0.00502574666958,0.000980911468344559,0.00481056290278925,0.00993791938207722,-0.0065386171265891,0.00888022757835838
"1821",0.00492987211074447,0.0062959344686595,0.0107046855690616,0.00791693673443739,-0.00563691688971479,-0.00352651971893614,0.00658285211667309,0.00983989511755623,-0.000240773745590395,0.000382775466384988
"1822",0.00819442760878686,0.00688197900710774,0,0.00662724017948402,-0.00246853871296671,0.0000978494260766016,0.00579682914442636,0.00292373052095174,-0.00762682253736069,-0.000765021771425012
"1823",0.00663076788160932,0.00683533661945801,0.00264783935353763,0.0117044323635678,-0.00854652000205469,-0.00206827894012485,0.00635450719156583,0.0021858199282192,-0.00177980744454487,-0.0122512563764504
"1824",0.00334656200662509,0.000411262927559219,0.00880299999772749,0.00192832216321759,-0.00574657276723478,-0.00434185947968535,0.000146670737785071,0.00799763150168586,0.00753708572442724,-0.00232554975998711
"1825",-0.00132369752149109,-0.00267323906349826,-0.00523572442126941,-0.00384911176026126,0.00438176746298957,0.000693745382226885,-0.00352363287201318,-0.00384700721842424,-0.00321751930501923,0.00815851687320612
"1826",-0.0118219061134838,-0.00371133677618907,-0.00438595952380005,-0.00265633413739375,0.00668277689006103,0.00614087784028827,0.00397807017551854,-0.000723990888735204,0.0133150583168988,0.00462429368806183
"1827",-0.0110515243597503,-0.00393207713491872,-0.0096916518707334,0.00435820754362815,0.00599257671477726,0.00236279283287399,0.0010273275446433,0.00458917724772911,-0.00525600063709475,-0.00230146453460378
"1828",0.00412286520771876,0.00332440386453148,-0.0213523263834662,0.0115720348688495,0.00238318162885354,0.00137482895321828,0.00557106793333007,0.00264479093214542,0.00944673734859536,0.0115339861699637
"1829",0.0107508308114288,0.0132532586991225,0.0145455469638154,0.00762637293761292,-0.00493752349007792,-0.000293808995460831,-0.00072885445317239,0.011511392751838,0.00182412568242118,0.00266054900521828
"1830",-0.0210060105132701,-0.018393604400786,-0.0286737440150915,-0.0106434729064873,0.00928033092329827,0.00421851414802155,-0.00890004099806507,-0.0113803886286649,0.0054623337555415,0.000379147925316126
"1831",-0.00900825359268143,-0.00666265015781287,-0.00369009766495809,0,0.00810276367841523,0.00205111668762248,-0.00603556355139456,-0.00167823320589511,-0.000629887400521389,-0.00454719271475734
"1832",0.00787804676159976,0.00482099358022214,0.0138887688122635,-0.00215145287923191,-0.0026188594969615,-0.00155956456224005,0.0037026282158128,0.00384337473988383,0.00724807374143221,0.00913592825592224
"1833",0.00688759521127835,-0.00438055371047363,-0.000913175702619395,-0.0150933261259981,0.00624749429763694,0.00117147576952981,0.0106239132482546,0,-0.0184591320838347,0.000754344303005805
"1834",0.0104779436245552,0.0111040547812804,0.019195598090386,0.0126490188148054,0.00125973264440282,-0.00155992088105483,0.00598621553624357,0.00885394428453035,0.000398462035197555,0.0018846720080643
"1835",0.00139679083002409,0.00580191175218037,0.00269041209727328,0.00912777077247795,-0.0109640970854885,-0.00566612137484224,-0.00275751305661998,0.00450644880032258,-0.00629282295449407,0.00225738301863121
"1836",0.00348734369755577,0.00185408994464376,0,-0.00618881376029634,-0.000817702339114823,-0.000196622843998462,0.00422078746515919,-0.00283350071217514,-0.00408819238476954,-0.00337844807662935
"1837",0.00454438416506875,0.0065804469083568,-0.0071556322063655,-0.00263470125504828,0.00336464379363455,-0.000392726913053365,0.00333308459835324,0.00497286115324536,-0.00370250327917743,-0.000376565178978328
"1838",-0.0023421450887664,-0.00326881138606694,0.00270280367172582,-0.00720491760512521,0.00571019012972385,0.00255561627971801,-0.00303311890156044,-0.00282745953076347,-0.000161552756192895,-0.000753569186683123
"1839",0.00202741423735531,0.00143484398068439,-0.0035939255906694,0.000967756434502975,0.00189277097702334,-0.000294306335619665,0.00333238768522337,0.00307181726233186,0.00646409168610051,0.00603313866066468
"1840",-0.00819880963439112,-0.00450260180942419,-0.0063117824454112,-0.0135332251246404,0.00143938032778257,0.00137302954184726,-0.00346582285578678,-0.00494712027207289,0.00698460191047867,-0.00412292080413723
"1841",0.00316708299226609,0.0032892520362382,0.00544437450685731,0.00489972215719536,-0.00485034635158632,-0.00146878024426977,0.00521667139409865,0.00378806438375223,-0.00438493980706378,-0.00338731004097692
"1842",0.00465537431349183,0.00840173543987377,0.00270780628703293,0.00950744717367891,-0.00135424027911324,0.000882769404397576,0.000576620124887794,0.00589611586169059,-0.000160121720694795,0.00264346846756669
"1843",0.00298286759540511,0.00792519476467546,-0.00270049387274618,-0.00193174381837424,0.00415778906651032,0.00264553203432039,0.00446629304522972,0.0014068166126886,-0.00512574078867745,-0.00527299793137248
"1844",0.000106011706019427,0.00201623411358387,0.0126354296611935,0.00120968358850515,0.0107278787979523,0.00287959194869436,0.00774516866277297,0,-0.00338108192415798,-0.00757290238187724
"1845",-0.00143365901603631,-0.00321938729147464,-0.00178252425720637,0.00555822474261514,0.00615959494416995,0.00146464466298823,-0.000426819652731836,-0.000234182438898944,0.010177665343029,0.00267073913185523
"1846",0.00191432156031368,-0.000201915783506923,-0.00267837708684493,-0.00552750164620031,-0.00603332246853483,-0.000584898273598422,0.00355955906622119,-0.00117093203289276,0.0092755718739097,-0.00228319130765142
"1847",-0.00870388998243488,-0.00222075107647723,-0.0026858896702826,0.00459170791732766,0.00401732866573057,0.00117065619464141,-0.00368898505139226,0.0042204816794631,-0.00190142606638066,0.000762844652970829
"1848",0.00588920059287945,0.0036421497653143,-0.00448839880881946,0.00529243927383494,-0.00355617981553191,0.0007795467612286,0.0116777486243769,0.00817164477723575,-0.0143673992451008,0.00266768573702603
"1849",-0.0010645586769692,0.000806686148989044,-0.00360664084886386,-0.00239314617251885,-0.00428296795788674,0.0010709190376188,0.000563117181499706,0.00115807300200088,0,-0.00304070567216974
"1850",0.0014918976241991,-0.00423063072143282,0.00814465104242279,-0.00167916334428819,-0.00322571618696343,-0.000778117159339176,-0.000140852389359458,0.0027756952785567,-0.000563743264294869,-0.00495612882897922
"1851",0.00973628823807426,0.00809228660531036,0.000897699483296099,0.0168190525559198,-0.00404529536710996,-0.00262853291725174,0.00211069816911724,0.00553643149486405,0.00676876723237352,0.00229889807629657
"1852",0.000895796068869359,-0.00220764431274112,0.0134527993805111,0.00378059999364488,0.00866486132261968,0.00390468680830725,-0.00589732632347217,0.00206468773342716,-0.00272133819879405,0.00458713250180853
"1853",-0.00473807038044072,-0.00140790958037917,-0.00530966526086762,0.00706223285339203,0.0108279538130009,0.00456899468130501,0.00254255636419098,0.00251861516179663,0.00971107559728845,0.00456614763446561
"1854",-0.00878010636554805,-0.00382667472187925,-0.00978649921415009,-0.00935039246432579,0.00796725445585245,0.0035808720171433,-0.00169081432071561,-0.00159921908166383,-0.00826644159075485,-0.0060605625859117
"1855",0.00346854260410079,0.00141521399323219,0.0017970121434645,0.0132138960811725,-0.00281023790378154,-0.00212199470768093,0.00733857871934762,0.00366011249583997,-0.00216395773416589,0.00114331630053921
"1856",0.00366924522719425,-0.00141321399301375,0.00179381331322204,0,-0.0073981774149956,-0.00125613058660801,-0.00364231546481708,-0.000227969231148206,0.000642586345381391,-0.000761353473580639
"1857",-0.00630510059351597,-0.00545899969633479,-0.0116385028428202,-0.00815101214936065,0.00221803865871584,0.00290273418812204,-0.00309361654573581,-0.00934555744964427,0.000882966754166548,0.00190477512353748
"1858",0.00842466041657564,0.00833502510654527,0.0117755526457637,0.00774842799040232,-0.00610895966638525,-0.00154361165684114,-0.00394915029836662,0.00437161758662619,-0.0024059908187346,0.00190111471928089
"1859",0.00243197954940855,-0.00100806893090311,0.00984763109133535,0.00698994006076648,-0.00142526416467392,-0.00106290686059618,-0.000849602948869377,0.000916339592161197,0.0022509767847172,0.000759081054928057
"1860",0.0040086091966729,-0.000403653733504261,0.00975179569051798,-0.00185113527248593,0.00535266869762463,0.00203099885102254,0.00751140634310676,0.00595111189676256,-0.0012833560805865,0.00227528168495428
"1861",0.00614663190727405,0.00868145739238257,0.00790169725768242,-0.00857672582347957,0.0058560128811016,0.000290131403774208,0.00604847254797924,0.00227516531803995,-0.0213637776666328,-0.00832387743504726
"1862",-0.000730995272185675,-0.00460351756999255,-0.00435539536238472,0.00584528504516912,0.012350087369396,0.00550054166213387,-0.00405490152017451,-0.0056752637780203,-0.0053344358692563,0.000381450015833007
"1863",0.00517285398483502,0.00361956622565396,0.0113734970373944,0.00278933292195349,-0.00531566240422265,-0.00124707561441062,0.0012636125330614,0.00525088498653803,-0.00214517332042496,0.000381422326485303
"1864",0.00161137279099099,0.00140262153968873,0.00173016833447481,-0.0136765568054023,-0.000437792393917058,-0.000769416392876199,0.00490727650205347,0.00272566421467624,-0.00421698355850864,-0.00762479245482162
"1865",0.00114208796638748,-0.00080036175319631,0.0120898332819503,0.00305531056989827,-0.00743363406248532,-0.00457549367760324,0.00181428135333728,0.00385069999430621,-0.00606163746574784,-0.00115257963929916
"1866",-0.000518514393954117,-0.0030036889722872,-0.00170636068428021,0.0056232684984252,-0.0123054167150216,-0.00503252140653287,-0.00125370129343927,-0.000677271108839639,0.00258984968896869,-0.000769141123897699
"1867",0.00202292638672597,-0.000803248259349187,0.00683732055956288,-0.00559182416972293,-0.000269144043685388,-0.000778212099512676,0.000976045101966694,-0.00293493965663116,-0.00208315970197215,-0.00269442259198116
"1868",0.00652180783798717,0.00824113086669098,0.00254680778650962,0.0105436150389238,0.000448300714366523,0.00145987001782522,0.015603424611202,0.00407613621920411,0.00751504663468516,0.00115791773421514
"1869",0.00478301383669355,0.00737644661897896,0,0.00996989064181419,0,-0.000777269393450242,-0.00205762846619995,0.00902085919784934,-0.00041441238473694,0.00424041755856797
"1870",0.0010235215547667,-0.00178116556712116,-0.00084667857998999,0.00367308491620455,-0.00143343924470263,-0.00145896295893622,-0.0107219232613455,-0.00446986257581172,0.000331655747187964,0.00422274939862954
"1871",0.000102248648403913,-0.000792991725915848,-0.00847447252848188,0.0052607348007736,-0.00367983418447393,-0.00175404422665215,-0.00514071423460127,-0.00202046633055641,0.00613341887884933,-0.00267588302880972
"1872",-0.00347640785939762,-0.00674607502962132,0.00256400987983052,-0.00341299778662352,0.00180183076033336,0.00136656518224343,-0.00405042224482333,-0.00517464835369341,0.000164799408228111,-0.00268298369309872
"1873",-0.00707974617206197,0.000199723010386732,0.00341011622002529,-0.00479452939901115,0.00890106316803663,0.00389815386143066,-0.00294478581687174,-0.00271361411541216,0.0101309196892869,0.0142198340612605
"1874",0.00304853047320575,-0.00139799643712102,0.00509754528258166,0.000458901626537944,-0.000534590135966462,-0.00194142712726952,0.00253130591242767,-0.00385494199079572,0.00260926290451113,0
"1875",0.000824087216171998,0.000199891064859958,0,-0.00458636070616925,0.0024965792120617,0,-0.00505048883059422,-0.00455277292416711,-0.00439168025692638,0.00303140980953276
"1876",0.00277918726033888,0.000200018176093941,-0.00169058724820492,0.000230507637030586,-0.00791623795129448,-0.00418257427275126,0.00112829741547893,0.00114319700888088,-0.00114359583636003,0.00113334305133139
"1877",0.00733971220519702,0.00799674098325931,0.0135477641614032,0.011054864396834,0.00771066460464431,0.00527451362934928,0.00619722147978319,0.00776624016028915,0.00318939322202638,0.00415104216286699
"1878",0.0011210836617741,0.00238020317477372,0.0175439409543112,-0.0056945132873365,-0.0128119036762194,-0.00252608385216613,0.0076985081401626,0.00317334635307409,0.0348088698917237,0.00977074474588324
"1879",0.0020301896631334,-0.00257228293582024,0.000820890814442032,-0.00206206102419138,0.0075704707592863,0.00116860928559914,0.00347284596104025,0.00246980795244167,-0.00346622020692899,0.00186078579704874
"1880",-0.000306281114880957,-0.00178540564831142,-0.00820334653608379,-0.00206600690595715,-0.00313063123949586,-0.000680971107952177,-0.00235314656315178,-0.00547550460502622,0.00276678260869567,-0.0037147358734172
"1881",-0.00602390192441127,-0.00765393439722661,0,-0.000460273574217851,0.0101391743526207,0.00408902503374731,0.000461805173536556,-0.00183545289020648,0.00102487191209888,0.00149140393515124
"1882",0.00451968584196027,-0.00123382358825175,0.00349772104339041,0.00211110690924854,0.0025761178441015,0.000969909827096327,0,0.00666536984571864,0.0000787131813189124,0.00148918296182177
"1883",-0.000715883957088659,-0.00144146643328091,-0.00331949705915224,0.00115724464375511,0.00478394411012806,0.00261529187040299,-0.00111894488273589,0.00616438226098182,-0.00204736596657007,-0.00408908711055656
"1884",0.0019441308023822,0.00123732279764788,-0.00249796571444472,0.00231202379856321,-0.00149861320513445,0,0.00602068156768731,0.00476487477352383,-0.000552347497379868,-0.00186641921430597
"1885",-0.000510344996804468,0.00041196315535208,0.00500844234615272,-0.00276801834172646,0.0024724766250237,0.000773197250559576,-0.00083503962621323,-0.000903198793715143,0.0108952230887345,-0.00598361722093199
"1886",0.00669308825328629,0.00885311786498821,0.0174418048826614,0.00948407116817895,-0.00837245343910831,-0.00326921886237841,0.0025072466847178,0.00565100533645602,-0.00265538908612728,-0.00300977948909364
"1887",0.0010149477439938,0.00102041404391984,-0.00244887013351025,0.00595771776692477,-0.0106874549382284,-0.00407582889364533,-0.00111150137182014,0,0,-0.00188676673158761
"1888",0.00491820897049,0.00550449090975391,-0.00327338408746769,0.00592271784440102,-0.00360123289807923,-0.00204634172839924,-0.0047295767833041,-0.00134867449694132,-0.0042286062074065,-0.00189041117318534
"1889",-0.00348121262675749,-0.0115571887087924,-0.00738923503891764,-0.000679144503998086,0.00731854466634618,0.00244131803070657,0.000978429214068655,-0.00472623736274702,-0.00110103016354102,-0.00795447621105305
"1890",-0.00643021405217936,-0.0133332208187137,-0.00330849196901972,-0.00453235231769167,0.0112117926207265,0.00457722004803762,0.00307172458926597,-0.00904560460340009,0.000393662424665209,-0.00267273931650935
"1891",0.00448439465324735,0.00395001069562029,0.00663897148264359,0.00569100265782074,0.000798162121290025,0.000194156153287661,0.00222716209616536,0.00890006576914537,0.00605962068151422,-0.00689125536772417
"1892",-0.00395695998074996,-0.0124249090370212,-0.0173124622299176,-0.00543251941109013,0.0002661583460839,0.00213242197953023,0.00319466319885531,0.00067822856566635,0.00547557119760866,0.00154199887714679
"1893",0.00137511359514941,-0.000629027368806767,0.00167788421560022,-0.00113775567874774,0.00637923151248754,0.00164459366838643,0.000692160003664011,-0.000451825706383913,0.00186716985428803,-0.00885304054897218
"1894",0.00503537661930764,0.00692404635446286,0.0117253555425232,0.00774682806027505,-0.00431392249077422,-0.00222112751390757,0.00456541200581695,0.00407039313681401,-0.02376143829602,0.00388352215418641
"1895",-0.00187260624573915,-0.00416755900240107,0.00331123053982019,-0.000678556874326164,-0.00203364537021233,-0.000870958297020774,-0.000275269783906684,-0.000450439181223117,-0.00946549467494828,-0.00928428552675742
"1896",0.00370152691517922,0.0079513642783684,0.00165003871410008,0.00248881584433658,0.00531606538592122,0.00145274708893695,0.00371937124856658,0.00743574691490889,0.00353330124093221,0.00156178810632168
"1897",-0.0113659338514825,-0.0153621369460677,-0.00658975411046026,-0.0187318171084634,0.0126038665237223,0.00580422317551443,-0.00590168973514926,-0.00849924478662123,0.0169640312317834,0.00233922971859379
"1898",0.010219018923237,0.0078010540833946,0.00497521900899245,0.0156394965073616,-0.00322088301421775,-0.00201961208249057,0.0088360122745168,0.00924858479076351,-0.00755369447017684,-0.00661216291621969
"1899",-0.00187130511501954,-0.00460267278852278,-0.00165019624858609,0.00339677581567344,0.00497748292073563,0.000288766085117853,-0.00287389207614086,-0.00223493112643014,0.00166494097355763,0.00469848805988504
"1900",0.00435784904724268,0.00483385536418135,0.00330568999992309,0.00925290896180875,0.00208551285303904,0.00125242961797767,0.00425460981462988,0.00403212743459269,-0.00474907407785574,-0.00428688944394529
"1901",0.00222011132487432,0.00104610422793527,0.00082382879459475,0.000894465773663811,-0.00130085519185752,-0.0000958886022791594,0.00218699821653301,0.00401602446861382,-0.000954310497126021,0.00273980957205633
"1902",0.0000502622693183685,0.00522350119538406,-0.00493829782357291,0.0044681800235864,-0.00746647033095471,-0.00404170671457904,-0.00259113469159877,-0.00177761448893532,-0.010109894679751,-0.00117094414663099
"1903",-0.00468156375704609,-0.00706715897677701,0.00330851452979086,-0.00400349648938014,0.0118087056748568,0.00386480036719239,-0.00560550219486555,-0.00823677959424629,0.011580241440776,0.00390772288067054
"1904",0.000404527339035843,-0.00167475924423599,0.00577092567972093,0.00692263799401638,-0.00138334407446272,-0.00115498496042876,0.00604938331591542,0.00157119880598899,-0.00166944111877387,-0.0019462560111887
"1905",-0.00429723925962688,-0.00293552603491976,-0.00245924165292732,-0.00598801913096558,0.00363667245756583,0.00134910696935164,-0.00464638808137718,-0.00112042550793923,-0.00302599931476344,-0.00312016237850077
"1906",0.000152358057204038,-0.0021029636909321,0.000821887677263433,-0.00490847213123313,-0.0138879609426051,-0.007024881946467,-0.000961165519798857,-0.000224360533350842,-0.00295523170020529,-0.00430358089483418
"1907",-0.0197480734653181,-0.0195996497209355,-0.0147784700778351,-0.0174886950420472,-0.00297403192742196,-0.000290703236434209,-0.0144314211736958,-0.0130162526585944,-0.0115357123842711,-0.0051080660694437
"1908",-0.00305568723336336,-0.0079536287255414,-0.000833076446691505,0.00547696893553695,0.00774076669275825,0.00588550892560424,-0.00195209909558147,-0.00250116582994531,0.0080233244835346,-0.00789890821798944
"1909",0.00722062978441862,0.00476693025359176,0.0016679060663003,0.00930569419662985,-0.00261850219207549,0.000579421776907951,0.00600813241046905,0.00364677294003046,-0.0031355443753549,0.00756371398691158
"1910",-0.0096961704714551,-0.011645133159359,-0.0158201315701111,-0.0152914239205459,0.00323802163312448,0.000482370983330371,-0.00888845949882666,-0.00885728762609772,-0.000967779675260627,-0.00474118489242559
"1911",0.000312729992388405,-0.00218226794395138,-0.0050762381848547,-0.00685084962680671,0.000610577328125306,0.000868178293522703,0.00182129119829,-0.00779094614222609,0.0145313228094457,0.00635168079479187
"1912",-0.00541468864517314,-0.0113710968333004,-0.00340123968372119,-0.00390884412209436,0.00932902097936417,0.0045296937785444,0.00153874109832275,-0.00461900805186355,0.00405826377111906,0.00197235968110299
"1913",0.0115687303813186,0.00906896666684753,0.0017064237982003,0.00900261482141018,-0.0021595723857526,-0.000864080792158495,0.00754183739688341,0.00556858677730743,0.0000792677127912089,-0.00472426408615978
"1914",0.00289777283441817,0.00197260600031601,0.00936959838756724,0.0128119544500525,-0.0000866541861963555,-0.000479716432763455,0.00554495493670615,0.0108442135665434,-0.00182267213213938,0.00158217528215698
"1915",-0.00139313069399394,-0.000437380893853034,-0.00168770376994021,0.00112909476556955,-0.00649323174443472,-0.00144146840369652,-0.00289509198591464,-0.000684758180719891,0.00023816291075085,-0.00631915096339819
"1916",0.00676900766944333,0.00415846271630604,0.00845324577846118,0.00541528309531736,0.00653566936019545,0.00327139549558386,0.01244320123776,0.0079947179698785,0.00166679104161904,-0.000794901731337117
"1917",0.00472168970282283,0.00566698473985761,0.00167622598274431,0.00157090375237012,0.00805098393200865,0.00201336534619667,-0.00027344182646194,0.00702443280314147,0.000871640274286101,-0.011933134359741
"1918",-0.000204029720230592,-0.00130041769420364,0.00167367202697766,-0.00268873229909639,0.0109068460114157,0.00401914129073,0.000956042733623486,0.00360036147608689,-0.00657109502923114,0.00402575128422056
"1919",0.00837926856469529,0.00781228760815122,0.00334175105868728,0.0096607390205754,-0.00993937469551331,-0.00314481590181748,0.00927978195564116,0.0047087946478912,-0.00414411848555662,-0.00842021728674447
"1920",0.00521896095765872,0.00193815117449025,0.0008327460823494,0.00467291229562505,-0.00308929994181517,-0.00105211924332282,0.000811233374854892,0.00490955538570659,-0.00224070904481988,0.00202189146360765
"1921",0.00267130281080252,-0.00429822713240768,-0.00582382774150259,-0.00199333676599356,-0.00163514864710812,-0.00296699264578937,0.00486337196618836,-0.00621807055907431,-0.00368943695861412,0.00282482003879458
"1922",0.00291593379387933,0.00561179104950815,0.00502101608093297,-0.00421684855678151,0.0056041028316518,0.00211165257256707,-0.00094107013688749,0.00335205147222872,-0.0107873449461653,0.00241449533829319
"1923",-0.00155387220207481,-0.0051514298842148,-0.00749380629913232,-0.00267414907226882,0.00557257638778386,0.0000961820892004805,-0.00672861987252471,-0.00178199131090251,0.00252282721002994,-0.00160580016755862
"1924",0.00507041895966953,0.0101404129110128,0.00335585996131105,0.00737427459102014,0.00375148499301181,0.000766092561214293,-0.000406499266948135,0.00401602446861382,-0.00365292631458847,0.00160838290910359
"1925",0.000649398298971038,0.00170864165123286,-0.00501693094176303,0.00598934644011062,-0.00322767936597823,-0.000191451247099073,0,-0.0013331810549605,0.00496985505898406,0.000401439712543361
"1926",-0.000399507351431572,0.00405137459954186,-0.00420166901916208,0.00507174794738541,0.00852131805400802,0.00277607288130555,0.00162647536068694,0.00311515729477119,-0.000243194166894112,0.00160511449347278
"1927",-0.00054925823666907,-0.00594625195512721,-0.00253153263721062,-0.00987278233255318,0.00523869332184512,0.00133675779769704,-0.000946933611286505,-0.00510185467177693,0.00551410963347387,0.000801271114856617
"1928",0.00284810073525588,-0.000213725141077425,-0.00169198709048135,-0.00155108799133163,0.00067245455540732,0.0000951494199421532,0.00501137256104456,-0.00267572775876646,-0.00112902419354843,0.00200165638693472
"1929",-0.000498255433916572,-0.000854686019717943,0.0101693597294445,-0.00155367384194083,-0.0172504745703967,-0.00638839553302739,0.000538858021850386,-0.00268266655261828,-0.0178427174403138,-0.0143828316073027
"1930",-0.000548272509536374,0.00940976242690339,0.000839102285492999,0.0131142630852707,0.0055684986671114,0.00144147042137899,0.000269606202886408,0.0100872928510416,0.00411015200805331,0.00405353459188329
"1931",-0.00144643576963543,-0.00508475586135282,-0.00335304641240308,-0.00263279173491859,-0.0121828314552003,-0.00355071921111549,-0.00188531371219969,-0.00754521822580179,-0.00548505107678998,-0.00403716978450852
"1932",0.00449529753481182,0.00212958337661906,-0.00420529424557281,0.00857884833716338,-0.00189736169397314,0.000288937102616238,0.0094444072788149,0.00178883385018058,0.00477440719193911,-0.0016213804612808
"1933",-0.00258560649560935,-0.0131748600930298,-0.000844518537007954,-0.0117773519964512,0.000432094576702458,-0.00105915503272447,-0.00173755917617435,-0.011160404945016,-0.0108962397328566,-0.00487208260272087
"1934",-0.00633114078615959,-0.000645683379021711,-0.00845308438217474,-0.0123593581622674,-0.000777256104475654,-0.00231311829767133,-0.00535569222026233,-0.00835232644653228,0.00115961232933959,-0.00815990734283745
"1935",0.0037628268706118,0.00409374800621021,0.0110827414644985,-0.00424585745595807,-0.00631007750755141,-0.00251213523966465,-0.0138643061415225,0.000455380442692555,-0.0050467525842619,-0.00699312305008326
"1936",0.00114932934614465,-0.00450638426465755,-0.00252955883876593,-0.00673239009688542,-0.00330538586840534,-0.00125931723960016,0.00122835130894328,-0.00750883103704703,-0.00656910848878922,-0.0049708498179174
"1937",-0.00584128820393837,-0.000646729906933152,-0.00338113691509812,-0.0106191708776778,-0.0104732507978463,-0.00378156015845144,-0.0287662521155861,-0.00320967204221045,-0.00912366276786081,-0.00791018072039307
"1938",-0.000753181760045685,0.000431423935869146,0.000848192432591155,-0.00502402893316722,0.00150001666134747,0.00184950404536055,-0.00407100299089669,-0.00850947910969291,0.00219633389583551,0.00125898658360835
"1939",0.0075384191237553,0.00366535919728372,0.00169485476286035,0.0130823872157899,-0.0040516076645597,-0.000291405294052804,0.00747050174952135,-0.00139172250765363,0.00160150877951359,0.00922045596687138
"1940",0.00134654444589244,-0.00386689228864101,-0.00846021236581751,-0.00928862354370485,-0.00256446005180389,-0.00252702417132378,-0.000699576956186054,-0.00627174432129363,-0.0108558527163871,-0.00415285260395082
"1941",0.00533021703985415,0.00927325161544856,0.00597271602382254,0.00137211221486,0.00319167879699167,-0.000682293657858102,-0.00727998600450641,0.00467499574226404,0.0020418410580072,-0.00959132395730922
"1942",-0.000901093145761922,-0.00491444461337853,0.00169629232584478,-0.00753604339975078,0.0127251757699567,0.00380285871686104,0.000563859351380147,-0.00503681648477594,-0.00585840555152328,-0.00294732818754173
"1943",-0.00772308989320758,-0.00365038000524232,-0.000846663704109685,-0.0151862199254711,0.00122207472776226,0.00213679640976161,-0.00887908766758094,-0.00329641778747403,-0.00204968834399821,-0.00844604763001489
"1944",-0.00572423858624027,-0.0129311841059101,-0.00169513214559902,-0.00560749437254637,0.00618808190500308,0.00213240211171573,-0.00568830957352973,-0.0068509200578063,0.00641848534734257,0
"1945",0.00782800964323616,0.00458520024430364,0.00594231895339914,0.0143325213403391,-0.00554402296578604,-0.00280505688122934,-0.00101041679060832,0.00404367372990677,-0.00467682831083038,0.00425901741067269
"1946",-0.0161356088019119,-0.0163007987438362,-0.00253153263721062,-0.0217743572428911,0.0118459236093744,0.0048499904126893,-0.00491196726912757,-0.0156363443306194,0.00290470731555637,-0.00212041208275215
"1947",0.00794546635238147,0.00419797135623634,0.00761419574445932,0.00449900713817653,-0.00146360611133944,-0.00212387340459785,0.0110339197627507,0.00890506342711306,-0.00281115088858641,-0.0016999779678657
"1948",-0.00181915080440453,-0.00748077142131354,-0.00587752525454943,-0.0202730901268559,0.00801749114844963,0.00319247768998188,-0.000287217155097053,-0.0102577223011575,-0.000256270293119143,0.00595994531177846
"1949",-0.00263225387493549,-0.00066479761142757,-0.00591202139044567,0,-0.00564475986145119,-0.000867653185884332,-0.00603275167361361,-0.00192796304902865,-0.00700675046575028,-0.017350806458111
"1950",-0.013552062331486,-0.0126444037218683,-0.0161428092882443,-0.0204524584507573,0.0193913551237979,0.00840181779842797,0.000577893506036986,-0.00748634589013175,0.00481884523551201,-0.0034453030602557
"1951",0.000154545758904501,-0.0112332875762298,-0.0189983744650919,0.0054041322478029,-0.00871199853430904,-0.00297247175606319,-0.00158849563241414,-0.00656921515043529,-0.000256906746345154,-0.00388940490539325
"1952",0.0110092428446804,-0.00431709853715223,0.0123241789061004,0.00855111973629796,0.00426626133409957,-0.000288863988159749,0.00679857968689812,-0.000734717702115195,-0.0182456487621321,-0.00954442786635024
"1953",-0.00117033330448824,0.00821528186163212,-0.00260900574230316,0.01308149273586,0.0005947180954331,0.00163549112371397,0.00129301933090908,0.00171542762842947,0.0123898262595776,0.0127025911314935
"1954",-0.0154362745303372,-0.0212764866125663,-0.00610273246082693,-0.00884764106489955,0.0135009643885806,0.00585841111971774,-0.00588298734985515,-0.00831880505153892,0.00284410930659407,-0.00389276939652727
"1955",0.0174892467523686,0.0191950398663752,0.00614020448606012,0.0149577119382334,0.000251417915135388,0.00353228151079632,0.0190531338247735,0.0148039746995245,0.00953936052303739,-0.00390789288984161
"1956",-0.019833106872155,-0.0297254980282756,-0.0252832379605511,-0.0156878957724658,-0.00435569141788694,-0.00171221038739289,-0.00127503167685883,-0.0133722760808217,0.00144716096495134,-0.011769807888793
"1957",-0.0114142420485447,-0.0137981096663137,-0.0143110060777361,-0.0217341413494089,0.0099267891090864,0.00390718106809906,-0.00141802188284124,-0.00566810618309155,-0.000425051006673338,-0.00352893522585584
"1958",-0.0164270748878809,-0.000236828188782345,-0.00907460538890459,0.0101209552165373,0.00608083259864611,0.00522119370894925,-0.00170419806021671,-0.00322160716818154,0.0079088445585116,0
"1959",0.00154749415930011,0.000711534914274559,0.00641020325195552,0.00586523369943781,0.00654093739102879,0.00198296384806618,0.0150803907260162,0.00273483411602449,0.00059060919483489,-0.0150509295657192
"1960",-0.0067663762084671,-0.0106659857711567,-0.00545933956403621,-0.0126337861023198,0.00789714276985976,0.00565526636232283,-0.00700786265088893,-0.0022316780009155,0.00337298265867214,-0.0125843292251807
"1961",-0.000858325529981552,-0.0103018829051812,-0.00365962155578181,-0.00910420412140578,-0.00636628121879623,-0.00271833054873216,0.00268188674279068,0.00447304106997271,0.00193296078549388,0.0100137531760711
"1962",0.0118109873172674,0.0220284878889256,0.00459135451983972,0.0111744963115283,-0.00558521166629211,-0.00291305226476601,0.0050675619293794,0.00890677153478703,-0.00192923165635606,0.00360527101475738
"1963",0.00970994633448696,0.00450013079759226,0.0201097192056179,0.00294710418686539,0.00363436414791396,0.00141399464652792,0.014285621833575,0.00882765123330298,0.00680733686540624,-0.00718459324177123
"1964",0.0198109112432707,0.0150908475423022,-0.00179224618526275,0.00416259004664599,-0.00798317352786371,-0.00272936232987786,0.00952776607366412,0.0109383390761726,0.00183634386052556,0.00814114085177753
"1965",-0.00711100627897532,-0.011149955581254,0.000897683080043787,-0.00658364323271299,0.00107869569644015,-0.000283168303021109,-0.000410319370843237,-0.00769411074943649,-0.00566573085316779,-0.011215776547182
"1966",0.0116248326015282,0.0136248742155722,0.00627797453578949,-0.000245580449958371,-0.00886716454337977,-0.00415371351123195,0.0075262198043542,0.0099345196957441,-0.00687111636906701,0.0117966179513764
"1967",0.00769485750961296,0.00463491294362317,0.0035652273161817,0.00712021217747627,0.00100322340311454,0.000852900077272345,0.000407471003053494,0.00239939158216385,-0.00143434866944858,-0.00627794142929505
"1968",-0.00137412179824814,-0.00553634279152482,0.0017760627992589,-0.00780111539328465,0.00183792647174763,0.00104193687509979,0.00597305335372456,0.00191483571483198,-0.00245035914576019,-0.00270768346460881
"1969",0.0114697735188325,0.0153097563504263,0.00531924977536002,0.0201472143446881,-0.00625325980090041,-0.0024601745322439,0.00323883046725837,0.0102720743675306,0.000338810779922261,0.0081448253341041
"1970",-0.00151187627637595,-0.0105095361723544,0.00529084048421535,0.00144517353271412,0.00226541296004634,-0.00331937469717303,-0.00739834688941499,-0.00638389168035269,-0.0143098562965259,0.0116697308327325
"1971",0.00641065436616572,0.00600307398344357,0.0078948152321956,0.00937945823641995,0.000836876287970245,0.00104672519244042,0.00853767999673982,0.00975688017762155,-0.0104802161161337,-0.00842948025412049
"1972",0.0114355248611253,0.011935117708721,0.0496082740816859,0.00428892711083684,-0.00259287115268114,-0.00161612358827534,0.00752496609298836,0.0254537228774463,-0.0219636943838234,-0.00134235562090357
"1973",0.000545405692432777,-0.0131552322999143,0.00663346702706846,-0.00830372165874615,0.000000220535217421158,-0.000371932255950558,0.00773539599748241,-0.000919395881731178,-0.00452691267435068,-0.00896049769793583
"1974",-0.00346933150217577,-0.0022981222564501,-0.0263590164418407,0.000956759943795182,0.00311000612550805,-0.0000951321190042487,0.00119102869851484,-0.00897199886879974,0.000624155138222893,-0.0144666273901938
"1975",0.00631619850593301,0.00691086307739908,-0.0050762381848547,-0.0088428988374325,-0.00142435049961331,0.000285836384733784,0,-0.00789189720459116,-0.0216538939435582,0.0027524450020886
"1976",0.00400303800184476,-0.00388930849727853,-0.0127550894972008,-0.0122981667551652,-0.00646190081634701,-0.00305250585021899,-0.00422976133662678,-0.0138044144000807,0.000819710348668234,0.000914806340723828
"1977",0.00093536409045436,0.000229696544334912,-0.00344511282456128,0.00634763965603535,0.0114873840322895,0.00641123634066432,-0.000796696216770476,-0.00450788880540942,0.0281216243571611,0.00457041564431049
"1978",0.00314761535285091,0.00459252902501706,0.00777853083338353,0.00266871698111237,-0.00918585598154509,-0.00408871576199354,0.00451710761010093,0.00762651844760542,-0.0222183055482137,-0.00955414996961046
"1979",0.000980532204672091,0.00731415709877647,0.0060034745286035,-0.000967832146026248,0.000674197490124318,0.000095514969519428,-0.00251293666886243,0.00614934451927662,0.0143038386230658,0.0050528032285897
"1980",-0.00107741909735071,-0.0115724808682206,-0.00511502379857653,-0.00193775931158802,-0.000842318370039785,-0.000381938664488435,-0.0051711295764163,-0.00376100189988759,-0.00481971612977761,-0.00319922509623971
"1981",0.00112764197156601,0.00367295036406845,0.00856897870913009,-0.00266917226066077,0.00236057970920833,0.00162347813227859,0.00399869672154862,0.00283147892060831,0.00152464573991029,-0.0183402430648723
"1982",0.000244777675041385,-0.000914897227430878,0,0.00827251485384539,0.00487748796918508,0.00209795335787089,-0.00610651386930194,0.0070587890827114,0.0250739057056308,0.0107426411771041
"1983",0.000636497651206103,0.00228939078665213,-0.0161428092882443,-0.0106178684055914,-0.0025107298224748,-0.00114192614044739,0.00373977877903453,-0.0042058050001792,-0.00366906609881124,-0.00415900323180507
"1984",0.00577387883048508,0.0139333795269143,0.0138169525022147,0.00536601939606496,0.00276873047400183,0.0011432316265263,0.00479041367763711,0.003754317850031,0.00876808394297024,-0.00510438663375412
"1985",-0.00160532203887043,0.000225402931300911,-0.00596247170117914,-0.000485056134431172,-0.00635885552549076,-0.00266436062712561,-0.00622465210293854,-0.00210365202113094,-0.0119078919102679,-0.00513052706809547
"1986",0.00175401432955979,-0.00427928264526023,-0.0102828071727715,-0.00169915367239226,0.00522036904197809,0.00181266909997735,0.00279850920104763,-0.0096042204303366,0.0103800228712174,0.00843884767950143
"1987",0.00535042611777925,0.00814281110142345,0.00779209560296468,0.0318502961058083,0.00603127730271535,0.00200007593660478,0.00730918623736088,0.00946054457357781,0.00461429562411375,0.0106925542322909
"1988",0.00280650033043428,0.00830153390517863,0.00171824579210078,-0.00824695380788465,0.00083256757573924,0.00114029688732398,0.00290250800138403,0.00163986542439964,-0.00242653611601129,-0.00873962635098224
"1989",-0.000723616606697508,0.00356055097155039,0.0025729477315386,-0.00641481865021021,0.00831951849145396,0.00246834874016577,0.00276219175574588,0.00233971106185882,0.00234554771657081,-0.00464030806755011
"1990",0.00255902446181056,0.00421265711627639,-0.00256634466086503,0.0126732029725345,0.00272303039778188,0.00170437439671822,0.00747754356157859,0.00210018412445367,-0.00190668231686641,-0.00233111440108369
"1991",-0.00211918242045783,-0.00684494091701304,-0.00343040983319887,-0.0200708331290741,0.00789929289216817,0.00387598561771196,0.00286441390996339,0.000465536405666711,-0.0264849157177869,-0.0457943004701402
"1992",-0.00694990824878694,-0.00111140509398056,0.00516342097096301,-0.0171083443732941,-0.00583416076522547,-0.00245272780054595,-0.00363543174450298,-0.000232473812891931,0.039871563287204,0.0205680919931677
"1993",0.00646393403408085,0.000222486954626788,0.00856154950503796,-0.000245168184261901,-0.00971197332273566,-0.00444443588014343,0.00351849327124154,0.00651918683738417,-0.0123520584602493,-0.0211132512505544
"1994",0.00386306759591371,-0.0017799134624652,-0.000848727395151183,0.0026974000931117,0.00390629781061502,0.000380097608283281,-0.000909110072426444,-0.000231484085430611,0.0103352701957204,-0.00588237341865872
"1995",-0.00110616491495108,-0.00401267154527041,-0.00254890121521767,0.00171192476020909,0.00836181028985927,0.00351286087337788,0.00155979769758607,-0.0115686226396319,-0.00386834859677898,-0.00295853949162506
"1996",0.00163695140679532,0.00492376536078987,0.000851897838427984,-0.00195326051061595,-0.00582942464707659,-0.00558194852127358,-0.00519080233876368,-0.00304291100505927,-0.012512918860362,-0.00247276535029672
"1997",-0.00668239930420345,-0.0075723037217138,-0.0161703782837974,-0.0146769862228523,0.0122221195485943,0.00332960220990697,0.00443537794663795,-0.0150269062023206,0.01179759678406,-0.0173525206683872
"1998",-0.000677875024605701,-0.00875217015864072,0.00519043372148431,-0.00943364527775714,0.00514030891435602,0.00369843676535386,0.00337662716671816,-0.00143013985929374,0.0208153655278578,0.0070634753146015
"1999",-0.0160312815760169,-0.0115463597796404,-0.0154904976458514,-0.0147873420213545,0.00730472589430931,0.00453541724308848,-0.00232976904554627,-0.00572970651021554,-0.00194604447168056,-0.0155310053935875
"2000",0.00507013011197865,-0.00366461783795857,0.00262206943970589,-0.00839478029956464,0.00411007364900273,-0.00169274447236478,0.00090800032258076,0.00432193196619024,-0.00228888608247602,-0.00916028487234122
"2001",-0.0161616084769024,-0.0236781479490337,-0.00959015762875437,-0.0164187684095958,0.0135622741384793,0.00819635106960503,-0.00907343676347661,-0.00812842635260913,-0.00237911458273243,-0.00821792272696698
"2002",-0.00686968543186184,-0.0174241424673961,-0.019366062631066,-0.014345270716338,-0.00205877454499437,-0.00364428204812084,-0.0117723022476712,-0.011086903418521,-0.0257218711959162,-0.0160538006646467
"2003",-0.00801950427086118,0.0119818576195743,0.000897683080043787,-0.00158769681022053,0.0123769301393815,0.00506442179186739,-0.00463273323776792,0.000974675263569091,0.00489551538504673,-0.00578939496770725
"2004",0.0196048913027389,0.0108925949826015,0.0167810092505662,0.0229868761841079,-0.00901251040782891,-0.00690540826620467,0.0223404365585251,0.00998325629533636,-0.00591561563938092,0.00582310723543245
"2005",0.0247288487341799,0.0210824267459637,0.0159715562718941,0.0136663449347862,-0.0177933839719331,-0.0056377345623152,0.00897510039304361,0.00867874275097202,0.00770110285379633,-0.00315774346202635
"2006",0.00425500501365184,-0.00145489773047092,0.00524015860263582,0.00700021654488769,0.0134459022542988,0.00368534609542692,0.00206265094539337,0.00320463810529259,-0.00330008678592986,0.014783378020544
"2007",0.00459996914192518,0.00439409343622565,-0.00260650369137883,0.0139031947052812,0.00135059900416645,0,0.0164671005983346,0.00816499333936349,-0.0193429821210155,-0.0182101106723288
"2008",0.00134953302730811,-0.00368411771420107,0.00174222595086215,-0.00914168820092831,-0.0198349168979481,-0.00828562986636472,-0.00506227646906521,-0.00119124493533562,0.0016880941353683,0.0100688091195851
"2009",0.0000962861706366169,0.00670225493450527,-0.00173919587866878,0.00230665789725082,0.00544272176529526,0.000722529206769629,-0.00411309236719182,0.00166968783844745,0.000266090123578033,-0.0131163498056155
"2010",0.00322462553958114,0.00114757910791696,0.00696869123317678,0.0079262412890484,0.00371146885950724,0.00133035231084633,0.00387197599245037,0.00428566532826102,0.0182673144879129,-0.00106324961847593
"2011",0.0013434171200517,-0.00802559290906424,-0.0103807556164052,-0.00608833118937402,0.00747518039812789,0.00341559350076515,0.00437114982628195,-0.00379337003472691,-0.010101924408222,-0.00957959621759008
"2012",-0.00536596738982698,-0.00970863966936053,-0.0122376320452308,0.00204190388804948,0.00271283283424362,0.0011357710729234,-0.00102429607489851,-0.00309386106374587,0.0134600072747426,-0.00107467628639846
"2013",-0.00992301912174109,-0.00723642468045649,-0.00530981444047729,0.000764071730331661,0.00190943625812623,0.00113248751230444,-0.015376709837104,-0.00763885361190875,-0.0140624569634321,-0.00753093793412274
"2014",-0.000535281421760514,-0.00493764159102039,0.00177954717979567,-0.013234718789659,0.0111180751212283,0.00509454495908868,0.0123633543243369,-0.00192435807647739,0.00440218340549059,-0.0119242345282613
"2015",-0.0180595458948037,-0.0300094745110773,-0.0115454375337561,-0.0177971678169465,0.0157084392509137,0.00610200487579915,0.00334276788489185,-0.00602561186082529,0.0150771473513824,-0.014262180473698
"2016",-0.00941901907685461,-0.0107186915624494,-0.0161724584748938,-0.00420200867257181,0.0180171320844809,0.00671773015001609,0.00730262951867466,-0.00339502272509262,0.01139896343526,-0.00946031160562877
"2017",0.0124611428197505,0.00935741754867925,0.0146118278230609,0.0216246857477227,-0.00197475084535292,-0.000185236296188274,0.012973682122692,0.0167884071744198,-0.00589141890646971,-0.00617957602536812
"2018",0.0177449638692677,0.0153694189426228,0.0126012224523444,0.0170365359545883,-0.0132429297780755,-0.0040789364757351,0.00565057842827321,0.0107683057354753,-0.00420852014085715,0.00395698354185292
"2019",-0.00801354400838028,-0.00624664408335973,-0.0106666351736541,-0.00329959107234123,0.0109525173912293,0.00493289822993837,0.000374546512618146,-0.000236838807395001,0.0113851990445886,-0.0016891660869599
"2020",-0.00783351768596374,0,-0.00359397710769649,-0.00814858394783557,0.00572187853416173,0.00351987184719205,0.0054919179704469,0.000947204076658048,0.0110864401997877,-0.0219966048061198
"2021",-0.00281270235059361,0.00435188256029839,0.0081155791555394,0.00872904070482861,0,0.000923028809454163,-0.00260712666309038,0.00828003629639218,-0.00337376861291772,-0.00403703159616031
"2022",-0.00603723400014489,-0.00192598066826988,-0.00178890329903403,-0.00559943657507245,0.00758645576453354,0.0046104699962155,0.00659617263253431,0.00375414645159267,-0.00160801450209835,0.0110017664138224
"2023",-0.0091604054007044,0.00603019941912497,0.0071683396517932,0.00230373477317025,0.0157354242520364,0.00853587365299635,0.00136021599661618,0.0018699291911537,0.0251759004392991,-0.0137458120305932
"2024",0.013114134304026,0.0141449878274191,0.00889677096943875,0.00842685093101969,-0.0127492385457777,-0.00737154442752419,0.00851949472888736,0.0177320964211729,0.0130642878606864,0.0191638030508074
"2025",0.00213254112314964,0.00732883347790247,0.00793675975594921,-0.00151952644154152,0.0132892402776372,0.00229181161603154,-0.0078352173855708,-0.00802377805364218,0.0137120473484831,-0.0136752043521947
"2026",0.00504807969444099,0.0077444153026458,0.00174968084698812,0.0220647638981257,-0.0115588774532464,-0.0047565998275283,-0.00148081628102259,0.00762655245959643,0.000241594208734153,0.00635480048784021
"2027",0.0148708470041266,0.00302752425783304,0.00436678699512938,0.0191065386203737,-0.00359781156619088,-0.00248167106781128,0.0195255633541802,0.00366973405970361,0.00804958525196198,-0.00114808995632198
"2028",-0.00548262731879212,-0.00510782963597789,-0.00347832102381385,-0.00754805693555527,0.0139177571249367,0.00654156846536158,-0.00206080363391614,-0.000228461252153145,-0.00798530684376009,-0.00632181185090264
"2029",0.00234177412959236,0.0151690626418217,0.0113437588895577,0.000490461746892379,-0.00304190229362811,-0.00228840858123602,0.00983841659636853,0.00617146454801309,-0.00998152596035917,-0.0034702855386991
"2030",-0.0131906128816066,0.00137957328158023,0.001725807630784,-0.00539462843048311,0.00156302322895896,0.00137650492001629,-0.00132279223979048,-0.00477039965199422,0.0114643794042504,0.00522343606937192
"2031",-0.0128242622209854,-0.0197429137632769,-0.001722834350116,-0.010847969600968,0.0163481682896263,0.00769649803452532,-0.00710593164505335,-0.00890229155914446,-0.00787784553251047,-0.0144341619889924
"2032",0.00924350118574035,0.0170959257994168,0.00862828952178196,0,-0.0065805729320173,-0.00354583533070585,0.00169834615585329,0.00967282218659826,-0.0215523905615361,-0.00468652079010523
"2033",-0.0125748545260406,-0.016117921963669,-0.0171087724435246,-0.0274178901285677,0.0177373501459435,0.00875994815346282,-0.0163480987867097,-0.0177915916204002,0.0222755461696662,0.0241318147701892
"2034",0.0123841271911942,0.0109993086848186,0.0104440220861803,0.0179395260554345,-0.0037754301462638,-0.00125046704455956,-0.00320076077959996,0.018810575718839,-0.00834345099255041,0.0137930332837239
"2035",0.0144610226652597,0.0217591199891845,-0.001722834350116,0.0188821230173251,-0.021166192537904,-0.00843722870188357,0.00926274381387349,0.00866198973170418,-0.0111909412055373,0.027777866916868
"2036",-0.00380786110984821,-0.0124601963479881,0.00517686141824858,-0.00494186361422544,0.00170901765859699,0.00164745767375374,-0.00293673843032161,-0.00949138938170757,0.00437834768166012,-0.0220628612013305
"2037",0.0100951586354994,0.0137644925479874,0.00858375901191244,0.00595971052168087,-0.0109793646580409,-0.00365403087754956,0.010431811758884,0.0182522324207859,0.00172724951920977,0.0135363096736323
"2038",-0.00276527047285513,-0.015388165107001,-0.00851070516971408,-0.0170327408617651,-0.0177016323581413,-0.0111845075639522,-0.0263570639330365,-0.0100828647922375,-0.0258642086717776,0.00278243448269144
"2039",-0.00447586004414968,-0.00390690668763249,-0.0094418579493305,-0.00150682120969514,-0.00160374264485752,-0.000463717907041583,-0.00474076730189488,-0.0140335906282935,0.00446728763037174,0.00998887909743806
"2040",0.0106532551602803,0.00945996239295699,0.0129982380264393,-0.0025151398247677,-0.00795392647381865,-0.00250401366492947,0.0035093559469066,0.00367322550884119,-0.00587393649196843,-0.0126373600584188
"2041",0.000580353601631112,-0.0061714303929048,0.0017107659101554,-0.00731211646461627,0.00185024957844382,-0.000371881011504316,-0.00212281531308334,-0.00251588682418213,-0.011817346063836,-0.00779065618397379
"2042",0.00961655834481667,0.0200091760730707,0.00683183985438274,0.0213361371581913,-0.00330892054432241,0.000372019358439557,0.0107645792990816,0.00985995564900533,0.00230627829503716,0.015142982519029
"2043",0.00411665463161071,0.00338216798446345,0.0118744104346229,0.0114397018457635,-0.0102685769302168,-0.00334774012937666,-0.00544884667310774,0.00681212251808616,0.00545429539643072,0.0110495723323076
"2044",0.00157290347452288,0.00247198781758584,-0.000838299991074765,-0.00221277357763516,-0.015055877604207,-0.00709072960892221,-0.00286402627512294,-0.00270644836346956,-0.0166977534319948,0.000546553163430996
"2045",0.0000951311456345305,0.00403493628874996,0.0176174775830362,-0.00024622218170256,0.00594012676665323,0.00479198557804406,0.00849143716378875,0.0024874693232193,0.00284453059487055,-0.0120152404922721
"2046",-0.000713749200333513,-0.00178602376478154,0.00741976644898523,-0.00419050194060056,-0.00661417215752902,-0.00252485825658733,-0.0190686788084447,-0.00383476723043108,-0.00343814692928124,-0.00331676100198663
"2047",0.00600055130656374,0.0134197906654152,0.00900153103821011,0.00668301693785045,0.00293284296075424,-0.000562817271106075,0.00921494044441151,0.0054348408424052,-0.00569262539774673,-0.00388247916964912
"2048",-0.000141805391118743,-0.00441404520628019,-0.0056771160479181,-0.0100809660031115,0.0114587303824041,0.00459702032259557,0.00787957941998996,-0.00180182100375326,0.00130118842211302,-0.00668153796059567
"2049",0.0028405383274972,0.00620696940876031,0.00489388260914092,0.0144062850738247,0.0131263350753521,0.00662987329274678,-0.0188631016612867,0.00518949662464285,-0.00147273672355541,0.000560530484758237
"2050",-0.000849751404133237,0.000660822878358447,-0.00243515663134941,-0.0019587982805821,0.00431840014808382,0.000927788057289103,0.00215012198916886,0.00246913257926162,0.00381741273959024,0.0151261328873129
"2051",-0.00118137798474427,-0.00462336620303561,0.00895050545415521,0.000245436661591603,-0.0136680434537548,-0.00593178913671655,-0.00845667705680275,-0.00335865745328245,0.00319795168188297,-0.00827820277748603
"2052",-0.0034059827081826,0.00176953376521083,-0.00403223478722536,-0.000735964721534255,0.00840782415335628,0.00354322562234732,0.00712889169396624,-0.0029204855566326,0.000775428620660046,0.0111296806566363
"2053",0.00631353505191479,0.00154556243316195,0.00242897764134797,-0.0014726841063768,-0.0186262640082127,-0.00744424877678374,0.00391798084482864,0.00856187959118038,-0.00413226569792469,-0.0143092756386252
"2054",-0.00410421950393092,-0.00859798237081355,-0.0048464249307113,-0.00762063971574189,-0.00362571442926107,-0.0021561545229607,-0.00264376226224061,-0.00513827768834441,-0.0018153440525589,0.00614179367706202
"2055",-0.00421556391174371,-0.00378014167592411,-0.00487004916024991,-0.0108990263800171,0.000316576187990636,0.000751535549684101,-0.00833176052150342,-0.00763538408257913,-0.00311769288024866,-0.00887895921922588
"2056",0.0010940949245335,0.00334829814943749,0.00570952971066463,-0.00150255818050582,-0.00126554617452634,0.000563381010428632,0.00331000506292645,-0.000452745533620513,-0.000955616358651601,-0.00391931914536592
"2057",-0.0140643989883698,-0.0180202306749787,-0.0016219671844836,-0.015299809276235,-0.0220916971771343,-0.0102269771853725,-0.0304490656485744,-0.0185643318080875,-0.0273043391304348,-0.0123666170244006
"2058",0.00414433635851919,0.00385143185130654,-0.00324929257765338,-0.00382055805893977,0.00923037763812373,0.00464491834478742,0.00889799296144766,-0.0129179718680199,0.000983372063442012,-0.00284572097699964
"2059",-0.0162215654116266,-0.0243735561314601,-0.01467005659221,-0.0222450628064117,0.0131576677307319,0.00424619489064781,-0.00492845580993129,-0.017060209566316,-0.0049120567570593,-0.0131278504276504
"2060",-0.00234174042346136,0.000693840974329785,0.00909832210480599,0.00758376028738184,0.00728564248025987,0.00178506304408788,0.00143386094431985,0.00285309753023166,-0.00601326523089696,0.00520530925471774
"2061",0.0127138849753912,0.00809052416241274,0.022131248810545,0.00622896433584397,-0.000707645892661479,0.00093814619091237,0.0165297470049208,0.0109054453212993,-0.000270871331828459,-0.00460298819676297
"2062",-0.006132452968026,-0.00710847078296961,0.00080191129730367,-0.0121228611083009,-0.00306823658312816,-0.0014992820577292,-0.00371298861074243,-0.00257961033783316,0.00144505056498345,-0.0202311155214705
"2063",0.0133606363073744,0.0145495878556592,0.00400649583883417,0.0120103981646256,0.00962756354096683,0.00347200025289496,0.0109240728533837,0.00940541309577125,-0.000631304129634969,-0.00118004618052503
"2064",-0.00297258103116305,-0.00409728934905795,0.00239423548439155,0.0116097593433102,0.00828509092282559,0.00205733202060543,-0.000890155960122208,-0.00652246752736174,-0.00541466483917807,-0.00708803408364778
"2065",0.0120216450241259,0.0237714287463384,0.0159236037298176,0.0244836451771657,0.0193026888536516,0.0114793635622084,0.0197225418499662,0.0192263102703472,0.0195989839361128,0.0273645963994336
"2066",-0.00456153737628451,-0.0136190820146114,-0.0117556082952225,-0.0169280595957948,-0.00509557221748846,-0.00470542054064238,-0.00149710141769621,-0.0025307204801549,-0.000711951569494884,-0.0167920756911898
"2067",0.00882706751408224,0.025124482865269,0.0158605308325934,0.0149405467650023,0.00527418985734585,0.00407839816016553,0.0242436445368563,0.0197230247559732,0.0113990470086467,0.0135453445761553
"2068",-0.00194858766319195,0.00507837852622051,0.00468365679263694,0.00299406502695465,-0.00121672429112896,0.00129294615109532,-0.00146384218185758,0.00136236523943389,0.00633971119133592,0.0116211714476675
"2069",-0.00561912248964136,-0.00175758432813622,-0.00233098494621631,0.00398021618310218,0.00966901524455976,0.00304277599069347,-0.0080647068200147,0.00702779309773538,0.00244989935733742,-0.00804142308010869
"2070",-0.0146537410673576,-0.00528150308551967,-0.00233628331142288,-0.0158574703657881,-0.00844530553649459,-0.00432090504455118,-0.0165175046884224,-0.00562799763857347,0.00139655232608882,0.00289521423429195
"2071",-0.00238155966198217,-0.00973466473343387,-0.0101486180233251,-0.00931524263361239,-0.0155890653036422,-0.00563150331458084,-0.00568247568020597,-0.00950852866613272,0.00653708690306587,0.0121247840176284
"2072",0.00228973622399264,0.00178732411210825,0.00394338829669594,0.00279552035761177,0.0124371563809789,0.00389993590411075,0.0034288370439135,0.00571394397544256,-0.00363703662182968,-0.0199657933908359
"2073",0.0122000246154679,0.00356845078907764,0.00392779256698828,0.019259944430815,-0.00495964517457737,-0.0000930289137738294,0.0112645269839133,-0.00454525009110462,-0.011385346973498,0.0052385780379427
"2074",-0.0087396407269531,-0.0162223137567461,-0.0195617449638658,-0.00223775325402276,0.00214710824499242,0.00259020670337673,-0.00725917334873272,-0.0109590823486659,-0.000791173626373598,-0.011580737745951
"2075",-0.00353614170746619,0.00880949559012811,0.00399031312850417,0.0124597238136683,0.0131344859163869,0.00475913898146385,-0.000126064268277215,0.00738706040815518,0.0170683963727469,0.0181605695309341
"2076",0.0035973455227909,0.00806094158694393,0.00874393633269754,0.0150134820614729,-0.0105953516507201,-0.00285119489357377,0.006682775387852,0.00801994599217704,-0.00276815748733827,-0.00517835431905656
"2077",0.00673325121302426,0.00932906707252212,0.0118203712783425,0.0128517209441479,-0.00558385100161207,0.00129132475201588,0.0100198888040213,0.0072744306571666,0.0122311156508599,0.0127241223596799
"2078",-0.00264668288914904,-0.00154038441243065,0.0046729678501618,-0.0050277470170762,0.00838432470242867,0.000828942202964811,-0.0162451449026906,0.00157980728080731,-0.0049704429690558,0.00513984965216796
"2079",0.00337720745904746,0.00110189934062377,0.00155029882825986,0.0209336990364595,0.00030548907386807,-0.00092013434814342,0.00277342573692074,0.00968912160612079,-0.00551201442156568,-0.0193180940344471
"2080",0.00442356838943314,0,0,0.00989850170284945,-0.0129643637206308,-0.00405388919919003,-0.0175990335117513,0.00290111453047692,-0.00692823238132634,0
"2081",0.00545700910343139,0.00330269491161306,0.00154798306794746,0.000700344466747715,0.00146783671607298,-0.000277104614484158,-0.000639880177308538,-0.000445079295315454,0.0113369061016291,0.0104287728250716
"2082",-0.00452280904592983,-0.0054860254841923,-0.00695508400084677,-0.00583049362825594,0.00138882358679093,0.00203501586828514,-0.0028167680722635,-0.0131344544515435,-0.0071570405522372,-0.00458721091733771
"2083",0.00191293910309054,0.00882616775625955,0.007003795990284,0.00445708496065711,0.00708778002897792,0.00295485503166448,0.00205423095539015,0.00902336299980955,-0.00607952932151745,0.00460835039256935
"2084",0.00448715478216322,0.0050304387207758,0.00463700205435447,0.00700605231275575,-0.000841309061598072,0.000552914062172061,-0.00589413178981091,0.00268280690022427,0.00865080376353022,0.0200688264583102
"2085",-0.000285113141849425,0.00174103648727386,0.00230752860982797,0.00788496062188293,-0.00497695780207996,0.000735788625910727,0.0041244566435843,0.00312160107545378,-0.00346531231049119,0.0106800103349713
"2086",-0.0115035236380383,-0.0134693184005579,-0.00767457416627282,-0.017487285969594,0.0114652938971305,0.00202267725397087,-0.00526289820721915,-0.0115585252542026,0.00495522042037044,-0.00222466379608099
"2087",0.00913685209903936,0.00110092859850752,0.00309365539145867,-0.000936802168555406,-0.008824888127831,-0.00183500952217219,0.00129042921779088,-0.000674675081100196,-0.00761243092755071,-0.00445924791956631
"2088",-0.00119137602677244,0.00769916797536174,0.0154200692910731,0.00586014321106743,-0.00452833086630844,-0.00211415508756463,0.000773373538296207,-0.00224999079232713,0.0057531031576612,-0.00727885080943291
"2089",0.00491435926085804,0,0.00759307434636614,0.0107203858125371,-0.0152660352556212,-0.0058042036928263,0.00296197452219205,0.00270640427080493,-0.0134338277023877,0.00338416449252255
"2090",0.00251608041455431,0.00545728394425815,-0.000753587447927417,0.00737835576581269,0.00430630752532868,0.00305767765114795,0.00179744059063558,0.00202415426386948,0.00729159259788115,0.01236644346353
"2091",0.00232073927933785,0.00434219608023589,0.00377073795453886,0.00366206759027055,0.00623713419687721,0.00351055616412554,0.00166638737232816,0.0060607871663545,-0.0140415222731023,-0.000555353763433186
"2092",-0.00415812332839172,0.00713364159583807,-0.00225386632966174,0.00387684713195724,0,-0.00156467770647051,-0.00268712100048163,0.00178496611146817,0.0201680578460488,0
"2093",0.00317883698307653,0.000429218016660515,0.00301195723624259,0.00159013609525371,-0.0137910061771865,-0.00461013090148665,-0.000256592689231172,0.00289529909297448,0.0086707706811624,0.00166675834314023
"2094",-0.00411452519542599,-0.00836729975292516,-0.00900890062575699,-0.0124745004412555,-0.0122555002440907,-0.00370492719731463,-0.0196354357917802,-0.00644025332906872,-0.00704891245510331,0.00665542577805445
"2095",-0.0100203704865912,-0.00302897772813437,-0.0257577218186668,-0.0151582691432078,0.00174947889252453,-0.000279299068814187,-0.0116508874667087,-0.00916408883409592,-0.0176608169394716,0.00771362090786609
"2096",0.0108412738013182,0.00802949442495038,0.0124418748294668,0.00606337848240956,-0.0134613879635896,-0.0054668176600714,0.00529787857505348,0.0024811753113283,-0.00343702297138437,-0.0010934787598561
"2097",0.0028472961103756,-0.00172239476049219,0.00460819713843152,0.0057950171816985,-0.00943518122976439,-0.00206013694895057,0.00263527043471257,0.00607599739097653,0.0090201271839383,-0.000547337882276788
"2098",-0.0114517316642343,-0.0148802219399641,-0.0191130812392187,-0.0108320408742525,-0.00138429151223962,-0.00168942029990404,-0.0219450351341258,-0.0136435125952145,0.00280455745494401,0.00821473346996493
"2099",-0.00411680640780543,0.00678644927041216,-0.000779410230338451,-0.0123484900106433,-0.0171206447665684,-0.00488835917972374,-0.00268696448389838,-0.00680272718209185,-0.000524357638950534,0
"2100",0.00398975438273275,-0.00413152139034834,0.00155988831780851,-0.00141546636965351,0.0134373799172745,0.0042512577722722,0.0132024215318112,-0.00639286818472562,-0.00821968338387813,-0.0157523714176044
"2101",0.0131659339837022,0.024890911388797,0.0233645013751749,0.012756832060153,0.00270121859278794,0.0038564794452709,0.015290197696612,0.0238971692833099,0.00484925947538795,0.00551868825165203
"2102",-0.00477271099637566,-0.00447384949530361,-0.0159816979883729,-0.00956373500641206,-0.0243247091265549,-0.0098389591621838,-0.0145364214030563,-0.0089767875856881,-0.00386068260190675,-0.00439071958871129
"2103",-0.00299134057044304,-0.0038517847726014,0,-0.00329730129810679,0.00259351174125921,0.000757025272519085,0.00292344988914128,-0.00181155444509351,0.00854400606486383,0.01047394718828
"2104",0.000190481026827172,0.00644467064314336,0.00618714302101031,0.00189050733921015,-0.0080107482135896,-0.00132375051951561,-0.00834734627587452,0.0111162627844086,0.0179039563318777,0.00109120500779669
"2105",0.010427743293679,0.0164353307568916,0.00538053340948474,0.00990561105712007,0.00269162016345215,0.00340877775410364,0.01817206160844,0.00964781631211498,0.00540537952624498,0.00599463697079994
"2106",0.00108381183815887,-0.00146984266137973,0.00458707979572326,0.0077067829123596,0.0200506571427748,0.00717182559436824,0.00826784567941252,0.00866633191238342,0.00298684929168802,-0.000541704379498187
"2107",0.0031065809319013,-0.00546800683090543,0.00837151497176469,-0.0101971494510703,-0.0167777205416891,-0.00674593132889489,-0.00299371157125272,-0.00837142243947475,-0.0000851016768919077,-0.00271010147902528
"2108",-0.000328269312835139,-0.00338330770521023,0.00075462255427583,0.00163909210715674,-0.00886669493808834,-0.0044338494021543,-0.00130542248605381,-0.000889008016197179,-0.0138699629136307,-0.0211955866319149
"2109",-0.000704359229199314,0.00297037068408623,0,-0.000701281173385859,0.00168798738162623,0.00217925383086803,-0.00209156842369551,-0.000444665277231637,0.00163951161998011,-0.00222107217221601
"2110",0.00291266661318779,0.00571189427984109,0.00377073795453886,-0.00350876192432548,0.0139859427700608,0.00595661404558911,-0.00458489164051645,0.000222372957620287,-0.00335975183735771,0.0122427460883201
"2111",-0.00238897618787692,-0.0094656106981601,-0.00225386632966174,0.00328628106035844,0.000415477252114993,-0.00225541132913332,0.000263067257722627,-0.00556028455535995,-0.000777975611064519,-0.010995183959485
"2112",-0.0107515793021554,-0.0205988827420454,-0.0128012368139586,-0.0159100791406158,0.0171094440914334,0.00621687783005553,-0.00605165676614328,-0.0138671970142267,-0.014619325512445,-0.0194552740661222
"2113",0.00949218857724343,0.012575898331286,0.00686504000384036,0.000237584735121033,0.0022867239726263,-0.00056137863722272,0.00754483352693369,0.00249471093566278,-0.000175621098213563,-0.0136053739085655
"2114",-0.00112828639852336,0.00064228581169834,-0.00227287428307532,-0.0130733876055154,-0.00244423949866768,0.000936496253675534,-0.000657054466851492,-0.00610842229110597,0.00114143472773232,0.00517234311863457
"2115",-0.00621289760722188,-0.0113416352799512,-0.0091115903927883,-0.00963385817036455,0.00220525068115274,0.000561178710976939,-0.0107796240768533,-0.0102437136876208,0.000701640081607779,0.0125786219037087
"2116",0.00203640912595904,-0.00692643524608527,0.00459777055074828,-0.00389113768139526,-0.0107476380272721,-0.00441211479321402,0.0097013689022063,0.00184012825446511,-0.000876406676185937,-0.00225858023963132
"2117",-0.000992724145909563,0.0076286112337911,-0.00228833287973562,0.00390633777952543,-0.0139520499531753,-0.00696271485791189,-0.00816028764330545,-0.00114785817077512,0.00403507894736843,0.0118846210882944
"2118",0.00264959872757142,0.0086523320742502,0.00382262868569572,-0.0051070060142564,-0.0160751072885034,-0.00852767304273749,-0.0120752069908314,-0.00459673931695181,-0.00716407484854154,-0.0128636462591393
"2119",-0.00844653704645837,-0.0113660564118058,-0.006854521053545,-0.0151552914977839,0.0130192229918591,0.00487403594357483,-0.000940734601908244,-0.00923599462112323,-0.00703980118831227,-0.00906514926579005
"2120",-0.00171313161748954,-0.0140997859321327,-0.00613509612626495,-0.00446750892255421,-0.0121798684356665,-0.00722802561333058,-0.012099438800715,-0.0146815146275207,-0.0053172458460562,0.00457409782496465
"2121",-0.00614959827986439,-0.000439983915517028,-0.00540114552153914,-0.000249330415946214,-0.00110539050543856,0.00143685762236379,-0.00204144735786183,-0.00402121881524042,0.00294014616785709,0.000569144195399662
"2122",-0.000143850426415515,-0.00506272835546406,-0.0100852123687302,-0.00598486453006397,-0.00791693976124164,-0.00325230506988039,-0.00722768374184135,0.00522458769519529,0.00222084036599446,0.015927265450697
"2123",0.0119930794711971,0.025000134727625,0.0164576178674962,0.01455073923432,-0.00875212100962774,-0.00383862811133617,0.00714270289735297,0.018190487546178,0.00850912072327614,0.0039193191453657
"2124",0.00322373040213719,0.00215810858299492,0.00462596225174328,-0.00494561234091917,0.0210349853691236,0.00789987766771461,0.00791044348213465,0.00255186151524223,-0.00457019691132188,-0.00892358463847098
"2125",-0.00765499017773719,-0.00969190554299504,-0.00537227474894364,0,0,-0.000573798194111741,-0.00189418039773015,-0.00485955689798001,-0.000264868439610377,-0.010129466925154
"2126",-0.00428550630649704,-0.010874289796337,0.0030866408515231,-0.0111829550693209,0.00161114779327654,0.00239137303936832,-0.00515189920410553,-0.000697739367321648,0.00441579075114928,-0.00454797665417239
"2127",0.00545168657038309,0.00065961669279524,-0.00461559950994483,0.000251419932364216,0.00787166838768671,0.00381661035317937,0.00844913159235916,0.00023240509703859,-0.00360505573889769,0.00285547202898218
"2128",0.00161711133801568,-0.00131836377083994,-0.00850059070470233,0.00603031365049445,-0.00772650007391829,0.000569860759040308,0.00621627343240916,-0.00302439389344311,0.00467700317684439,0.00284745874768899
"2129",0.01039936172247,0.0127612099694838,0.000779262294557048,0.00924065356865778,-0.0049089458082261,-0.000759888793650632,0.0138329252351521,0.00560090237887323,0.0129117437489985,0
"2130",-0.00443928364462243,-0.00391048611150291,0.000778887807170614,-0.00866133601621433,0.0128433687368259,0.00532358996501903,-0.00649097435944956,-0.00359041387731085,-0.00173427852930974,-0.00908585572589227
"2131",0.00512317215619462,0.0233370562562201,0.0155641552067913,0.0144782371381589,-0.0204064250302567,-0.00841606328323352,-0.00986660106439863,0.0101273336279182,-0.0128561845155615,0.00343846653051139
"2132",0.000708033508354022,-0.00149186957653658,0.0114943744333482,0.00984276822675856,-0.00600067097152934,-0.00305176420338871,-0.00484807960157541,0.00373020506989108,-0.00659978886483448,0.0119930413004823
"2133",-0.00726285208881006,-0.00787786230800114,-0.010606109874057,-0.0070664575880921,0.00862402553679531,0.00296566909518581,-0.00562477957789642,-0.00766529639524172,-0.00265748075699779,-0.00677197507159488
"2134",-0.00304031042886987,0,0.00200097246859188,-0.00343618807021773,-0.00350554421112603,-0.00248015338424523,-0.00947437873324453,0.000702219598581078,-0.00133221427594676,0.00113634815293406
"2135",-0.00019078219574975,0,0.00460821940299394,-0.00942719890863131,-0.011241023084764,-0.004780493507058,0.00485177131175951,0.000233665257202142,0.00106720026561358,0.00454040856141935
"2136",-0.0209700632810045,-0.0335599562343512,-0.0252293793219545,-0.0222889887433528,0.026468847370684,0.0116248636537495,-0.0160022537456919,-0.0240877542906661,0.00453093469315813,-0.00451988643037415
"2137",0.00209296594641817,-0.00748970449930952,0.00470597495388425,0.0148566199005866,-0.00693262268324002,-0.00275427792785343,-0.000420609382057124,0.00311514269782576,-0.00619082869019183,0.0215664003574805
"2138",0.00801571978275128,0.00548814370178352,0.00702564601085265,-0.000757168457274915,-0.0134976743444498,-0.00522623499194463,0.015287437575612,0.00334469312237617,-0.00347067713435945,-0.0122220558958132
"2139",-0.000915722723323964,-0.0002275189398252,0,0.00479907129402646,0.00328607341917153,0.0035470615644102,0.00221047884115078,-0.00214289698402959,-0.00196464541977193,-0.00168738161556348
"2140",-0.0028458418621915,-0.0245677463598537,-0.00697663067339305,-0.0279034200011654,0.0185347988918061,0.00707016856308784,0.00454836194509833,-0.00978276378239684,0.00268428771144791,-0.0326760730635546
"2141",0.00628864525023864,-0.000932681593462714,0.00234179776477283,-0.0149986837493136,0.00939494234143323,0.0026563864201492,0.0153678576341314,0.0019279487744619,-0.0116008925861304,-0.00582415211058229
"2142",-0.016777303951266,-0.014706065428325,-0.0412771615979164,-0.0343921973992904,0.00863654305569139,0.00397358260729286,-0.00527029757367659,-0.0264555451071835,0.00297936072626648,-0.00468652079010523
"2143",0.00180901211257778,0.0175313362515475,0.0121852131180118,0.0193040493718217,-0.0197022121980049,-0.00697350743554559,-0.00475476818413756,0.00963430061938886,0.00243050688380619,0.0117715903659563
"2144",0.0125915564494359,0.0419091522691211,0.0160512172206979,0.0253398085420107,-0.0158583839866886,-0.00692849071295132,0.00696164741866001,0.020063758519276,0.00116735810733348,0.00465380499809842
"2145",0.0110371461381868,0.000670533341460944,0.0134282716684846,0.00676401917808733,-0.0031022418738692,-0.00267537971376297,0.00149098835840111,0.0115136956257664,-0.00448470722907357,0.000579150118952709
"2146",0.00433811439280207,0.00848599470016631,0.00623529077560958,0.00180870689289936,0.00328445458376248,0.00316191516590392,0.00270680400022894,0.00758812774880524,-0.00225245521673045,-0.00347241290050826
"2147",-0.000332331978333711,-0.00465019110832954,-0.00077459466577845,-0.0113489999819608,0.0105972779094659,0.00382059462085116,0.000945048323354847,-0.002824083658437,-0.00523743914100483,-0.0116142449742631
"2148",0.00802441999871184,0.00912127424723441,0.00387591290059119,0.0125229096246389,0.00690551903959036,-0.000380602196395907,0.0071478374276146,0.00991274694006372,-0.00363110008601675,-0.00470034876032666
"2149",0.000847867447957951,-0.00352725277059718,0.00231666891479132,-0.00128833305720744,0.00516462317687671,0.0000955465236649466,-0.00388339702031582,0.000467380590163158,-0.0101129735766586,-0.0053127963211177
"2150",0.000517555345493914,0.00309728355771499,0,-0.00645000364314752,-0.00421166279148966,-0.00199878869884884,0.00174778930122543,-0.00186877066306257,-0.0271514491090392,-0.0160238240596492
"2151",-0.0039512183775311,-0.0037495277127978,-0.00308171091841491,0.000259731551730535,0.00541366276314559,0.00276518458564867,-0.00362332656918074,-0.00397852698626777,-0.00312198684357579,0.00422195857957752
"2152",-0.00179460435611178,-0.00730575441686443,-0.00463670988986586,-0.014278499929954,0.00622547582468691,0.00123705158273602,0.00282823882021122,-0.00258436301425735,-0.00540950919399696,-0.0144144029424824
"2153",-0.0056298719794815,-0.00289917244495264,-0.000776482597506956,-0.00974451885067695,0.0124584788020243,0.00408447088487907,-0.00711795123857506,-0.011072211393378,-0.0044847422380323,-0.00853139209343812
"2154",-0.0103719869764008,-0.0118540602973378,-0.00932394189529828,-0.0143614983129285,0.00247739076651765,0.000946252548491788,0.000270550180041518,-0.00262031736881474,0.00977663165385545,-0.00799018329028789
"2155",-0.00581749034740209,-0.00792233822888477,-0.0039215964243291,-0.0188885465042907,0.00535448585296661,0.00330822497491123,0.00216365604021762,-0.0028657778496558,-0.00465113440248954,-0.0192069322486307
"2156",0.0122832618781812,0.0134612263637814,0.00472458751465887,0.010176214688481,-0.00729199193095809,-0.00282658841723793,0.0018891076565164,0.0124551633177932,0.0015258058218024,0.00821227311896955
"2157",0.00687887309652235,0.00225132475439871,0.00391843791884727,0.00980117236630584,-0.00371477179788182,-0.0014169743518162,0.00511798020425625,0,0.0014283089343452,0.00313291822478545
"2158",0.000237213429243877,-0.000224708155990405,0.00156126168898196,-0.00997571723645219,0.007704880017533,0.00113545538699245,-0.00375206359455404,-0.00260243194116438,-0.00855758312365851,-0.00374779901424127
"2159",-0.00151780901476872,0.00629069855297137,0.0077941187262327,0.0108932015964092,0.00739972973925029,0.00585836663366646,0.006456126739256,0.00308358700171429,0.00632974987042534,-0.013793109233514
"2160",-0.00337300969095089,0.000223252488680048,-0.00386692012852963,-0.0167024781986888,0.0105263840083587,0.00304924892839686,0.00494441767143949,-0.00425615839996396,-0.00791005432192893,-0.0165288315302095
"2161",-0.00195418346960508,-0.00267853299718046,-0.00155286046872471,0.0035616282617299,-0.0079317574985347,-0.00515973113735668,-0.00518607172454666,0.00403688678512171,0.00201729110503912,0.00581769849731795
"2162",0.00329535619161359,0.00671436769818978,0.00622082966701987,0.000272849882013482,-0.00750614934488392,-0.0038658676640978,-0.0042775657056292,0.00496669252385251,-0.00364296814577625,-0.00385605447913029
"2163",-0.00818767447336977,-0.00111162278171673,-0.00309115382533776,-0.00873348050422051,0.00887754939073093,0.00350235715209579,0,-0.00117682411338627,0.00442604637736932,-0.00064521886644664
"2164",-0.00191996961715912,-0.0040063257456594,0.00310073868558702,-0.000550693664033597,0.013118560271244,0.00396163425243579,0.0034902185180774,-0.000942470341302903,0.00249068878715097,-0.0038734139922495
"2165",0.0125992539180155,0.0118437442743728,0.0146832621202542,0.0168044786335639,-0.0123851814611373,-0.00413416191818017,0.000134099770577434,0.00778317597879385,0.0102245482995786,0.0213869496870762
"2166",-0.00902322696486024,-0.0136925657757676,-0.0175172062151208,-0.0219454836760518,0.0158791228761086,0.00660503414174118,0.00668788512711549,-0.0142756740395733,0.00510784141971388,-0.0133249515791739
"2167",0.00119791439519035,-0.00582186648346783,-0.00620145645838888,-0.0155123178519413,-0.00545059294835104,-0.00037549550126581,0.00146183161504387,-0.00261182372725011,0.0140221905887035,-0.00321539024234307
"2168",-0.00124423297495413,-0.00292787753730828,0.00780011421873894,-0.00168812077928804,-0.00322414237231095,-0.0026249743492609,0.00199008315905869,0.0016665460349865,-0.0082598515081207,-0.00451613365891079
"2169",0.00364228175505832,0.00158122616145739,0,0.00140893753250326,0.00234503010455134,-0.00103431316682612,0.00569374146649992,0.00617868158810064,-0.0000936084587908059,-0.00648092618506435
"2170",0.00558678312386118,-0.00360839399780821,0.00232202740308063,-0.0109765315932372,0.00451740788950805,0.00178807628215583,0.00750512795138847,-0.000236051000548687,0.00262048671259696,-0.00391384098282155
"2171",-0.00289665816014018,-0.005658886248044,-0.00694977759190962,-0.010814060135763,-0.00787031215804435,-0.00159691402062678,0.000783930750768658,-0.00519717834764355,-0.000186651736768018,-0.00523909389894606
"2172",-0.00790541159711255,-0.00956068315264735,-0.0108863208058256,-0.0123703406666167,0.00987563929586233,0.00611585173602691,-0.0054846226075066,-0.00474961873262914,0.0134441414112207,-0.0111914887418054
"2173",-0.020881377319044,-0.0216042511988987,-0.0298743461908856,-0.0157296202873517,0.0100992922128704,0.0027119857249589,-0.00774647288948083,-0.0174182151402661,0.0174113214902445,0.00266307934858157
"2174",-0.0301024255058043,-0.021611324966379,-0.0340356933225653,-0.030778334802554,0.00301570495647896,0.00401077229206215,-0.0195847207361083,-0.0206412568681417,0.006247690940824,-0.0166002437314864
"2175",-0.0421068655336458,-0.0268907692789102,-0.0352348257364755,-0.0436640344914877,-0.000316674593418553,0.00167182149448086,-0.046699965814751,-0.0453755541663535,-0.00539906430484294,-0.0249831944517125
"2176",-0.0117678807987023,0.00616817270045433,0.00608687296800836,0.0127713028135317,-0.016065180205917,-0.00547139680851738,-0.0252018135139198,0.00701281332751114,-0.0123947798099592,0.00415521063827451
"2177",0.0383939215060984,0.0166747790970849,0.0397580652682827,0.0331021777847089,-0.0193037525634874,-0.0061547067708434,0.0249817766090461,0.020118668659816,-0.0136497429956122,-0.00620695348291322
"2178",0.0247351133912244,0.0108541181514457,0.0182876006150599,0.0442478364765475,0.000574290762656693,-0.000562772962100944,0.020121858372621,0.0199746921732753,0.000557304737759834,0.0360860590358638
"2179",0.0000501466132800665,-0.00238615697177935,0.00489805568691937,-0.0128580632065616,0.00295102697287142,0.00018762132162653,-0.00111115053323141,-0.0101634382988658,0.00900393551460321,0.0261219592799926
"2180",-0.00807915793508773,-0.00454442849140002,-0.0154347187023525,0.00177604208841475,-0.00768218557549905,-0.00168971234381488,-0.0198859806652854,-0.0120209239338691,0.00110398347113105,0.0241513737615482
"2181",-0.0298476406212245,-0.0285920857338701,-0.0453795722233137,-0.0387112607481843,0.0072050967141597,0.00449212352366923,-0.019012477418793,-0.0263627672389302,0.00349197757765118,-0.0331421357263799
"2182",0.0189811955092778,0.0140984930958568,0.018150584318078,0.0144479868310672,-0.00860410556567504,-0.002718688361521,0.0107031182919965,0.0179637770856582,-0.00531130051221518,0.00856963182897941
"2183",0.000716345607942204,0.00146344896062267,0.00763994257779532,0.0039394779177504,0.0048765515157978,0.00244392379879232,0.00200318857156567,-0.00306890142807303,-0.00718106222110859,0.00653585802039114
"2184",-0.0151367926079241,-0.0211883942115232,-0.0320135339286063,-0.0298823055565421,0.00913054176245964,0.00309485295083656,-0.0189944766303699,-0.0218057402262927,-0.00324553053581345,-0.012337627793219
"2185",0.025130944050316,0.0291116653825398,0.0234987124174919,0.0317360797201094,-0.0147539778904292,-0.0043939844409624,0.0151405370640112,0.0251770284089683,0.000279086431837161,0.00723212063576195
"2186",-0.0133716585604472,-0.00531920019536269,-0.00170056853691969,-0.00512651303208156,0.00479880979627523,0.000375728701073941,-0.0121899121141957,-0.0138144655264477,-0.0129278277416619,-0.0130548529148178
"2187",0.00544173944022575,0.00947979923058706,-0.000851767166973549,0.0103061956902502,-0.00675193846277766,-0.00225281826750412,0.00116152598342234,0.00985731479992991,0.00235560168724014,0.00859783403115144
"2188",0.00454422719902303,-0.000963027235667768,0.000852493292770262,0.00390040588815266,0.00630032120793023,0.00263395017452717,0.0163860553304584,0.00205505749123436,-0.00206799216209796,-0.00131145753062911
"2189",-0.00371066790794239,-0.0106050666656551,-0.00255541639653756,-0.00149452669328987,0.00156530861540793,0.000938411872074996,-0.000570661118391547,-0.00281984638556843,0.000565156346452156,-0.0124754099800847
"2190",0.012499558590636,0.00682103617884944,0.00768582072454271,0.00957801140366032,-0.0191644823081587,-0.00787409231791081,0.00842272051498094,0.00385612482018138,-0.00301260588389562,0.00332449124458023
"2191",0.00866648651116031,0.0164529582078587,0.00847436121075895,0.0243107063171968,-0.00377358472896949,-0.00028298631158441,0.0128820802438014,0.00717038059877217,0.0133144095691329,0.0165673099142225
"2192",-0.00224800577793816,0.00285652931903368,-0.000840246977840353,-0.00231530176439187,0.0122054419878075,0.00831662916734999,0.00978369106160804,0.00101692921942198,0.0102507317165359,-0.00651901687994838
"2193",-0.0163413352754319,-0.0256351051861363,-0.0319596169840316,-0.0185670411035254,0.0153844972287067,0.00468631930315011,-0.00332191299012363,-0.00787767676589268,0.00737934665144002,-0.0150917261893305
"2194",0.00516775383708845,-0.00219263747697684,0.00608167852039587,-0.00177348275588685,-0.016297928951256,-0.00569104236649143,0.00874848358988012,0.00438259581012823,-0.0062265360885132,0.0113257646300211
"2195",-0.0129795929787723,-0.0302732212309329,-0.0146804386689416,-0.0186557210214856,0.0139037073980735,0.00497303989514775,-0.0132155838832505,-0.0148869968938511,-0.00681837286297216,-0.0059289081563676
"2196",-0.00159883849822984,-0.00377658033853157,0,-0.0159926245091431,-0.0000816410985048366,-0.00112084808949275,0.00460381458970294,-0.00338703178676814,0.00398923829678788,-0.00795224601006539
"2197",-0.00361573033707863,-0.00404317130477838,-0.00701147604992203,-0.00429317914491001,0.00681611640478574,0.00149572600066628,-0.00916543322420749,0.00967290298017653,0.0209757621421571,0.00601201054571754
"2198",-0.000259308375677558,0.00659710919100509,0.0247132415039764,-0.00215587919062543,-0.00864610544236977,-0.00261305582978888,0.00503656261221641,0.0137238157300856,-0.00615440322480598,0.00597601393501157
"2199",-0.0250971276869755,-0.0186537512087048,-0.0241172266571912,-0.0212964531140641,0.0171136292047986,0.00570801210455296,-0.018018173186532,-0.0153258823588482,-0.0126582280786489,-0.0138613336739144
"2200",0.000585067393215066,0.00436661332499977,-0.0123565016986178,0.00473049436454565,0.00283140192223241,0.00344265248142084,0.0070243463003079,0.00337222968102879,-0.00405824578598513,0.00669341801839107
"2201",0.0186581454516572,0.0179028088553228,0.021447877400584,0.0288762107932132,-0.00346874570230704,0.000185553226346835,0.00996408363331769,0.0170633214866418,-0.010372309398806,0.00731379861976911
"2202",0.00260940677213095,0.000251584616074441,0.00699892326073082,0.0054913122237441,0.00426639990484734,0.000779369288711695,0.00465111354182435,0.00152508768251569,-0.00121652628470403,-0.00660057038275963
"2203",0.0149375890656682,0.0198438189875771,0.0121632632875579,0.0266988029233171,0.00605793041153757,0.0048242338606288,0.0086985135557458,0.0114211338585366,0.0211748799444895,0.00664442739342297
"2204",0.01779508409289,0.0189657321351868,0.024892794561189,0.0215722965557883,-0.0135676679025509,-0.00553953316725975,0.0179413059586313,0.0225847184935524,-0.00201854302263582,0.0132014125057576
"2205",-0.00342633315757668,0.00459278912865391,-0.00837517838415092,-0.00173564826746997,0.00431315387083719,0.00204253490309858,-0.00245941489826684,-0.00319017070086935,0.0100211825876946,0.0195439748149826
"2206",0.00819055102041144,0.00962449083946959,0.0160472556337674,0.026659051779975,-0.00332258658984219,-0.00250167076067098,0.0097247602801418,0,-0.0014564354500598,-0.00191690668555067
"2207",0.00902668543823326,0.00881808348021385,0.00332495917271536,0.0107253553344606,-0.00837408940916862,-0.00260089579917966,0.00827463112160243,0.00960101403589286,-0.00510481326631207,0.00448137263945814
"2208",0.000596253569710603,0.000944933704173589,0.00248555033317666,0.00363028584191949,0.00262348261921996,0.000559018079372198,-0.00107616856932158,-0.00414497409946968,0.015851237088613,0.00446151072916767
"2209",0.000943767143757546,-0.00354026975672717,0.0016528731041372,-0.00751286061466849,0.00760549891320261,0.00335059048826936,0.00538692390115636,-0.00195915486205489,0.00396856668254975,-0.0158629878376184
"2210",-0.0063021786613805,-0.0106583556531175,-0.0107260021949709,-0.0162598926227694,0.00170425817256881,0.000927705935070522,-0.00736758037612684,-0.00981354396547585,0.00494118237249452,-0.00644743147882887
"2211",-0.00479392346442531,0.00526687958461358,-0.0116763939386997,0.00769453199000036,0.00875046219566755,0.00546791802998636,-0.00647776536146027,0.00941534237547459,0.01743247794178,0.00259568152702783
"2212",0.0153543475777316,0.0126218523402915,0.0253163384090249,0.0243212107839732,-0.00489931532842558,-0.00341033248543265,0.0114100524286311,0.0130093146329633,-0.00456899226024055,-0.00258896140772769
"2213",0.00454676285628297,-0.00188147621264889,0.00493845800636539,0.000828244501405617,0.000322891963484784,-0.00083231388311833,0.00805789629717779,0.0031501627834265,-0.00706154994208186,0.000648920381757012
"2214",0.000491752421426073,-0.00376983223344773,-0.00491418948794387,-0.0102067559420689,-0.00274367778769757,-0.000463021768109195,0.0118570859031295,0.000966030408747764,-0.004178158132779,-0.0181582545830651
"2215",-0.00127834823133388,-0.00307471324471931,-0.00576121608773472,-0.000279017339173238,-0.0061491368709955,-0.00342659118488542,0.00118519781824222,-0.00120651304840635,0.0063382076326961,0.00198147886929001
"2216",-0.00620324647366366,-0.0045078781082698,0.0132450999617693,-0.014496641046729,0.00993226703160754,0.00343837308378481,-0.00355104527592343,-0.00507371347566343,-0.00887075289086969,-0.00856956398348829
"2217",0.016893707787156,0.0102478613577182,0.0122547233144297,0.0206507240412339,0.00169278990050059,0.00101875423233455,0.0109542406381198,0.0179698367895273,-0.000358014847632204,0.00332449124458023
"2218",0.0109612855253851,0.00825666184375184,0.00968533441098152,0.00582039252104161,-0.00853037978479798,-0.0056434691463394,-0.00913837331119527,0.00238561203021459,-0.0017011549520789,-0.00596420155884292
"2219",-0.00245746228271038,-0.00491359814382897,-0.000799254032444963,-0.00909357435704283,0.00665583324974461,0.00260478487641214,-0.000131468289243153,-0.00380787662244608,-0.000627802690582935,-0.00266663025528879
"2220",-0.00193243770462748,-0.00940477088083047,-0.008000055767866,-0.0114014830781868,0.00249955616991127,0.002506083714231,-0.00250364658579971,-0.000955414908062391,0.00224356097998735,-0.00467914912177814
"2221",0.0113747359115455,0.00735792700218063,0.00967736987739065,-0.0115331010191829,-0.00402152554393675,-0.00518382320473232,0.0038308578326387,0,-0.00805874820916908,0.0167897693851011
"2222",-0.000574328312508254,-0.00424116798418439,-0.0111822136101104,-0.00939085819740304,-0.0159089477137155,-0.00614138973976852,-0.00105265968151946,-0.00645656319695886,-0.00956849620480682,-0.00594450458779516
"2223",-0.00430967204187893,-0.000709961330592424,-0.00484644815128099,0.00172361788628517,0.00754973650033786,0.0019663715521967,-0.00724558011692478,-0.00216595590159729,-0.00382790736576821,0.00996670947658385
"2224",0.0118309996393469,0.0113663792181171,0.00730516348776766,0.0197876428670234,-0.00459525618281609,-0.00287319038484501,0.0221600813373226,0.00554749563566581,-0.00649594675674436,-0.00526308626300498
"2225",0.00289916976269011,-0.00210723110898059,-0.000805694481556984,0.0132171235855298,-0.00820027779846655,-0.00262788112455414,-0.00986613606407205,-0.00407776926187475,-0.0148263473552389,0.0178571708144006
"2226",-0.00303307391301266,-0.006804201831349,-0.00483880459692088,-0.008048851842135,0.00115764938371421,-0.00103474856263519,-0.00432653417853068,-0.0144506682901088,-0.00944103544285746,-0.0168941229624917
"2227",-0.000998477324019809,-0.00307094760198834,0.00729332381586012,0.00167876740509398,-0.00264274812525134,-0.000659634814402232,0.00289692047750667,0.00171077907114814,-0.00311410773696219,-0.0079312219733344
"2228",-0.000523428693689709,-0.00545048814594695,-0.00241338970956828,-0.0139664166095658,-0.0146559489970882,-0.00678684111643013,-0.0286239946346352,-0.0124421220526897,-0.0145778210391692,-0.0059960575746596
"2229",-0.00933122578356715,-0.010483752890379,-0.00403228640000508,-0.0249291585143203,-0.00563033717405981,-0.00170809504721026,-0.0135171914666325,-0.0249506174847026,0.00288188286036273,-0.00871308670317672
"2230",0.00230676131743901,-0.00433412696309399,0.010526333264772,-0.00435788534289416,0.00295768679619668,0.00190138828792175,0.00918078350923279,0,-0.00210729881020499,-0.00202843934733932
"2231",-0.00393177607946549,0.00507866115338063,0.00400643845496096,0.00204270857604927,-0.00210658404537156,-0.000474682557072947,0.00122178011061069,0.00810751525217102,-0.00335955077750061,-0.0101626021929274
"2232",-0.0139599123617533,-0.0153995994720076,-0.00957713827991991,-0.00961008227173354,0.00481327862698988,0.000569689088637748,-0.00718741715887306,-0.00804231208428485,0.000192584027880471,-0.0143737315317003
"2233",-0.011228280201404,-0.00855327246426307,-0.00483473209066154,-0.0138192641785628,0.00571418516771138,0.00379511756860529,-0.010517683509159,-0.00481388837512708,-0.00279248922084718,-0.00763885608064085
"2234",0.0152069542581563,0.0125708810217,0.00971663716545068,0.0193797933889139,-0.00091905729575914,0.00132329594070391,0.0117338084425771,0.0132385970434059,0.00144844537366651,0.00489846340708389
"2235",-0.000729478718535126,0.00316472304187387,0.00240582102855802,-0.0029246818209181,0.00167277870574578,-0.00028343163539768,0.000546087688451546,0.00477377832667147,-0.0132099413095164,-0.0153202689780357
"2236",0.0158659892265629,0.0101917185122535,0.00480000756232979,0.0108534064266399,0.00208720759777425,-0.000472115668945339,0.0106365448877097,0.00725168215289695,0.000879460655831998,0.00424322340568328
"2237",-0.000862207733270837,0.00576498979080142,0,0.00899620136762369,0.00666569383507354,0.00217291830222521,0.00283381121768067,0.00570978362088792,0.0110319047154153,0
"2238",0.00364397864102695,-0.00740380760371384,0.00477692720169642,0.0100659659796767,-0.00306251731103491,-0.00131944263651362,0.0102258438135845,0.00444347469103201,-0.00453845122708474,-0.00140843151233594
"2239",-0.00114668636956805,-0.00697804397786905,-0.00475421665483533,-0.00939639485606936,0.00307192513493892,0.00132118586547536,0.00173176557652033,-0.0105675124878224,-0.00805115949369128,0.0077574441065984
"2240",0.00133946748752822,-0.00169605908871551,0.00477692720169642,0.00517392250393045,-0.000082925460024974,0.000942700911534811,-0.00491953285030966,-0.000745118712761728,0.00664971627909816,0.0160951672652541
"2241",-0.000143406450846428,0.00582526897442115,-0.00633906954925956,-0.00772074575908976,0.00231783456506407,0.000564964812391766,0.00334010096050896,0.000248515249163805,-0.00466293948585716,-0.00137739162486072
"2242",0.00114670429256081,0.00482622180509673,-0.00478469681817928,-0.0219021702635001,-0.000990958229333705,0.0010348612200568,0.00799060523735529,-0.00472170925727278,-0.0118094769842814,-0.0151724188841127
"2243",-0.0041517908244636,0,-0.00801296337623991,0.00147319419476455,0.00396770046041484,0.000376645297502698,-0.00634151819116047,0.000499522708796496,0.00661726419753084,-0.00630257884926444
"2244",0.0095358505095815,0.00696452947990722,0.0153474489989149,0.00764937350870309,0.0135074862850624,0.00531805423094989,0.0123650991902249,0.0187168753378446,0.00353219198454058,0.0112756100009341
"2245",-0.0102049984020699,-0.0114477017006201,-0.00795539841506265,-0.0119710146468306,0.00032580026225193,-0.00280876227982385,-0.0189125806416606,-0.0142084695391501,-0.015545532025279,-0.0209059238447552
"2246",-0.0140028455779136,-0.00506619019628884,-0.0096231326768349,-0.00561445207104205,-0.0271834774663611,-0.0105165206069423,-0.0147255964147782,-0.0067098193542805,0.0106266757249642,0.0113878176129558
"2247",0.0195029167979159,0.00994161382070557,0.00566785085112587,0.00683496331493938,0.00878446162577506,0.00370086129218028,0.0167121423388858,0.00850648867434334,0.0222090699251363,-0.0014074403706511
"2248",-0.00605849834486072,-0.00672266513327857,-0.00241541990233729,-0.0165288649611878,0.00970324690836288,0.00321435504293643,-0.00267288318984538,-0.00868282487583816,-0.0129782641697249,-0.0288936282311872
"2249",-0.00671951960775918,-0.0157117065966428,-0.0129135542207369,-0.0111044217583951,0.000492588855885989,0.000565692220448444,-0.00241161482319041,-0.010260237494752,0.00165577094878278,-0.00507975678233286
"2250",-0.00777982262141064,-0.00221043425296319,-0.0114471699849166,-0.0081941668466905,-0.00106711628717138,0.00150683383719485,-0.00617870326634862,-0.00278142124138148,-0.00194473947665263,0.000729459707354385
"2251",0.00258138553488996,-0.00319955110916903,0.00909828687358782,-0.00673210969364346,0.00131510731200346,-0.00216306637437447,-0.0056764967415236,-0.00329570643345434,-0.000876812167544982,-0.00364433985582713
"2252",-0.0193812214244437,-0.0170368201626206,-0.0155737092468744,-0.0280345212523885,0.015758183896744,0.00801135048036072,-0.00462129895790742,-0.0167900162349679,0.00546073119081236,-0.0102415653600367
"2253",0.0050524799991174,-0.00150719389991216,0.00915898218077094,0.0161648871408626,-0.0129282534965196,-0.0073865211764832,0.00314057955369584,0.00491602061606899,-0.0128018619648738,-0.00665179463204035
"2254",0.0104979017142119,0.0090563579992069,-0.00412544196235187,0.0152838034807081,-0.00589403468984939,-0.00254360659332475,0.0110260910968747,0.00334718401401246,-0.00265255916443108,-0.00223211243083221
"2255",0.0146317892307775,0.0184494333269769,0.0248551010161888,0.0196622104050981,-0.0021408630465517,-0.00264423562054772,0.0196584599060967,0.0207849612031843,0.0121158691523602,-0.00447421180545382
"2256",-0.0152380261151588,-0.014198321074159,-0.00970092734747641,-0.012955930090176,0.0113054876201086,0.0041661527725072,-0.00488586163616367,-0.014579996765361,-0.0218978102189781,-0.0104869787599111
"2257",-0.017815142243892,-0.0124162175809316,-0.0122448969704209,-0.0033575307149285,0.00554851581446281,0.00358325533264381,-0.0127388710364092,-0.00282331093306309,0.015323393034826,0.00454210752137274
"2258",0.00824902924727033,0.00475441551094047,0.00316363501699124,0.00780741925835304,-0.000243124898365976,0.000470091591874278,0.0051072750665262,0.0036034695415994,0.0108780967181683,-0.00452157006397669
"2259",0.00907445249883065,0.0072992388403792,0.00746886830648608,0.00802459516454834,-0.00722389847567839,-0.00281743779342802,0.00414560066855962,0.00487285196021858,-0.00523510411565486,-0.0045420296094798
"2260",0.0123833915010487,0.0194902312538829,0.0107083907105192,0.0140844528320503,-0.00752224203110108,-0.00226024278627612,0.0113200553022379,0.00995445265305328,-0.00292372085641046,0.0182510150888562
"2261",-0.00165059399788148,0.00147060771321961,-0.0122251242683519,-0.00362315312971428,0.00572930357390899,0.00183403633835777,0.000266347658576693,0.00151642468596225,0.0072329685706769,0
"2262",-0.00228498311851155,-0.00416045169626511,0.000825159992828173,-0.00696953777337306,0.00295494727692613,0.000188312612783736,0.00293358027833968,-0.00656099701182888,-0.00756919919740318,-0.0141898071176862
"2263",0.010671976512129,0.0088471944516828,0.0148392430242072,0.000915337288331264,-0.0166136830905165,-0.00528328006886136,0.0102363907992755,0.0104140940647039,-0.000684462716861178,0.0166667524346811
"2264",-0.00708780948524623,-0.00803874107681501,-0.00568648873967359,-0.015548803104815,-0.000998300364370985,0.000379336673877351,-0.00447415676052942,-0.00703870989962796,-0.00763208437276164,-0.00968705542198245
"2265",-0.0100032829426557,-0.0149805357157816,-0.00980394495034864,-0.00309702224658992,0.0044981322776978,0.00113796952291878,-0.00753474030992607,-0.00962039310664209,0.000394409394486317,0.00526712378627625
"2266",-0.0139794694698046,-0.0149589773104761,-0.015676448895698,-0.0273375535366791,0.0072151996262777,0.00426157917774161,-0.00972292386560225,-0.00894687694481067,0.0140942244637712,-0.00748492787745059
"2267",0.00169131612468632,-0.00632735446862465,0.0125733339909304,0.00223579895328263,-0.00403459463954126,-0.000282983604974585,0.0164092858192764,0.00154784844093969,0.00281855382270924,-0.0098039421145949
"2268",-0.0126142977989183,-0.0168111397738384,-0.0173841182014508,-0.0191205480743303,0.0134755095777703,0.00603758333353976,-0.00330854304635564,-0.0100440095908986,0.0144407637138981,-0.0159939228439159
"2269",-0.0239916427499774,-0.0181346656092086,-0.015164280894201,-0.0308642939863112,0.0017947242214813,0.00215642228024882,-0.0223049386028144,-0.0228927994164445,0.0141397155658682,-0.00464405853976857
"2270",-0.0109764325804312,-0.0100263404236193,-0.0213858817272133,-0.0107274612447024,0.00447833959979471,0.0025260536729439,-0.0118140053464484,-0.0135783661037202,-0.0044277154135145,-0.00466564641415823
"2271",0.000989856518493371,0.00346493973090278,0.00699321883096804,-0.00033885562809266,-0.0109435178469989,-0.00317305925118661,0.00398521407356811,0.00377895422949681,-0.00889479560938689,-0.027343700059397
"2272",0.00806851690563226,0.00796802289133547,-0.00520851907234643,0.00203389704901502,0.0144253740181868,0.00449399909840809,-0.00698074460589448,0.00430213592721551,-0.00506013948940498,-0.00642569783124736
"2273",-0.0249405558789701,-0.0171276854501491,-0.00872605145266192,-0.0104871999582878,0.00985658532189748,0.00391452018642147,-0.0151619712424005,-0.0109774568822159,0.00489398334990865,-0.00565877484512667
"2274",0.0164165469432167,0.0128684998380684,0.0123240638616968,0.0129916076488972,-0.00936037713771132,-0.00204233908271922,-0.00139947689914854,0.00893348110084102,-0.0162338042758421,0.00243899091980437
"2275",-0.0214660033302023,-0.0367920092116133,-0.0278260423244094,-0.0394870889233299,0.0155870031668732,0.00465152139117975,-0.0113524601776094,-0.0300508687020815,0.0102893130544353,-0.0210869089061161
"2276",0.0013311824892579,0.00906849976457935,0.00805007766095378,0.0147574683883072,-0.00310159943540622,-0.00129620442400535,0.00297725727031151,0.00553238976276793,-0.000960789758632008,-0.00828489181420122
"2277",-0.0128151226685028,-0.0206971352927823,-0.0381544767233861,-0.0218142790489818,0.0105296796218639,0.00491407748197226,-0.02657295501708,-0.0220080508160693,0.0133679549903456,-0.0075187801837816
"2278",0.00560208471160628,0.0108454800856879,-0.00369001265020841,0.00389389298329634,-0.00678867782500847,-0.00249124276281953,0.00667954903294365,0.00450067539958332,0.0011387965890064,0.0134680023834841
"2279",0.0205152131238875,0.0264097236004661,0.045370486459378,0.0342030641873465,-0.00381496648211377,-0.00221982906283202,0.027693529423144,0.0229626636397564,-0.00464497117537155,0.0299002652026497
"2280",-0.0151165413483058,-0.0134011998189386,-0.0212578685755503,-0.0170474664264765,0.0054253190679614,0.00333718671441341,-0.00982434014658073,-0.00848620562336033,0.0102857333333333,-0.021774146157322
"2281",0.0136430260711764,0.0214614921821286,0.0135747711780834,0.0145680729481956,0.000476238067402157,0.000739356613040476,0.0214031198571365,0.0168416330434895,0.0114064760292898,0.0197856396611851
"2282",-0.010883144675219,-0.00851066186933813,0.000892821275057187,-0.00341867693316134,-0.000238133034898502,0.000738189107056808,-0.0155424511428918,-0.00705951935132443,0.00372822253958227,0.0121261125018888
"2283",0.00520920716502937,0.00214619298378405,0.00178407360311206,0.015780460119674,0.00142817221180835,0.00129173162990215,-0.00662577294771205,0.00710971049011166,-0.0106788093475939,0.0111821204449172
"2284",0.0243772867420784,0.016059835732168,0.0240427565844004,0.0324214934055871,0.00847634506365291,0.00534410159017051,0.0217118058795283,0.0285096175137194,0.00384828229915257,0.00947862482423667
"2285",-0.000361521902392581,-0.00158072100487816,-0.00608685215063798,-0.00948639397707429,-0.0030614516447004,-0.00230359869084695,0.000138750037508295,0.00712774546915895,0.0102852363801376,-0.0187792482003014
"2286",-0.0180221038364191,-0.0274404043199921,-0.0104986872950545,-0.0323646210806806,0.0185523134947561,0.00708360817716702,-0.0105541620875704,-0.0212322040358289,0.000370134186854276,-0.0175439474833902
"2287",0.00599505789537247,0.0151927582462399,-0.0123783783732585,0.0283276370550229,-0.00829335779086071,-0.00109600834515045,0.00491225940009055,0.0182108790606041,0.010731834979437,0.0251624127265246
"2288",0.00156812134788575,0.00133591532674249,-0.00268604094276359,0.0076336307121172,0.00484564673266386,0.00237753969422627,0.0011175754361803,0.00236726877202109,0.0120823798627001,-0.00158359108553852
"2289",-0.0190501585216495,-0.0152120250867369,-0.0170554542308498,-0.0115284740484218,0.00116647841425221,0.00127730187146091,-0.0224611964314704,-0.0170559116299508,0.0158270778692231,-0.00634416643820135
"2290",-0.0134609473461123,-0.023577436866375,-0.00182650845372834,-0.0136620800523344,0.0215199933672963,0.00747153482604856,-0.0293989861796693,-0.0149490343650436,0.01344375,-0.00478852442938482
"2291",0.0000541011086510057,-0.00888154296209476,-0.0192131872350615,-0.0138512809369771,0.00106426188550102,0.00018081320582497,-0.0161740362969401,-0.00406516525137612,-0.00219625753850028,-0.0256615684840983
"2292",-0.000863110311586479,0.00420060730190452,-0.0177238685485288,0.00411099399176229,0.00881294887615236,0.00298413288371568,0.00523095253853989,0.00027188639107889,0.00774781638056332,0.0016460680853132
"2293",-0.0130080152623532,-0.0142218954632493,-0.0199431346465897,-0.0167178567560625,0.00700328622524782,0.00459764335861235,-0.0147192703887982,-0.00843283037533582,0.0401887038283129,0.0123253916243458
"2294",0.0206170398057774,0.0195191760306186,0.00872104814303509,0.0173490258013167,-0.0166018302228368,-0.00762787062202286,0.0129772525665279,0.0150893451081413,-0.00587936344497497,0.0146104412805887
"2295",0.016878094142398,0.01609287759583,0.0365033111683206,0.0221691283476813,-0.0105702214629541,-0.00298417700262155,0.0192165445519819,0.0202701256871944,-0.0303312265095367,-0.0112000939303752
"2296",0.0163348064844782,0.0207540261821471,0.00834097017973834,0.0196863164980472,-0.00614878917261852,-0.00244916380410742,0.00906161714631204,0.012715016239053,0.00618633805488367,0.0210357295389787
"2297",-0.00409598634460817,-0.005885727790782,0,-0.00589001314610849,0.0122961907393506,0.00463739329659241,0.00955965693934258,-0.00392367428611728,0.0243331999220679,-0.00554667519181595
"2298",-0.000468426915899989,-0.00188369527600141,-0.00459562583676154,-0.00460830405041557,0.000840061161214489,0,0.00215218712856258,0.00787839530880774,-0.00600218948345443,-0.00876506550734024
"2299",0.0144794811842524,0.00727976252123419,0.0166206995279345,0.0248016443555237,-0.000534085051709488,-0.000995859510952601,0.0115962323021692,0.0104220133099917,-0.0177751655421812,0.015273351601643
"2300",-0.0126299719073619,-0.017398499411745,-0.0163489682392385,-0.0212971783698916,0.0040475634858963,0.00199310556682053,-0.00240582424856439,-0.0167612696400335,0.0149796781536007,-0.0134600760332335
"2301",0.00457569587817996,-0.00435832869427955,0.0101571092680075,-0.00230796837442904,-0.00197800784746838,0,0.000425396651227317,0.00550738826323771,0.00332707726218162,0.0128411642829631
"2302",0.0121118570001946,0.0139534098620515,0.0118828885929345,0.00330478680411628,0.00358237312346743,0.00298385357763431,0.0181511816068918,0.00834639154134531,0.00263580475609393,-0.000792463724620274
"2303",-0.00230121462538357,-0.00296803188275385,-0.000903233641757706,-0.0098815234669124,-0.00964455273288711,-0.00486779373961321,-0.00306425902413876,-0.00646666601726287,-0.00686903844757536,-0.00158593958574915
"2304",-0.00784260743137699,-0.00460107016341793,-0.0153707423103369,0.00864941075439241,0.00437094331514176,0.00163048266288324,-0.00167643529707284,-0.00104134741521478,0.0130646228924549,0.012708406021543
"2305",0.0235069378687986,0.0274607439212458,0.0247934028600945,0.03562002794313,-0.0176087397045241,-0.00781611344013522,0.0260286815828188,0.0242376379996825,-0.00733312548325293,0.00078430302575816
"2306",0.00449259552195125,0.00238177767880354,0.0143369185948776,0.0133758567998801,0.00412704081663318,-0.0017344083823605,0.00763764490494867,0.0058526378045114,0.00772695103320764,0.00548589929572096
"2307",0.00391945208929623,0.00844751246289599,0.0070670673356219,0.0113135622245235,0.00364417412620122,0.00118871018922984,0.00500817416712573,0.00455345511472549,0.0172733653522075,0.00545596840250417
"2308",0.00325349979234479,0.00523570069372581,0.0105265052121097,0.0198881728255198,-0.00641251871475657,-0.00337925263262073,0.00269354380635689,0.00302173650660942,-0.00157377615570831,0.0193798199127144
"2309",0.000798348902588897,0,-0.0104168521635167,-0.0015233381174814,-0.000311192146765449,-0.00201598407063375,0.00188028667424001,-0.00577433987422071,0.00497758416311944,0.0182510150888562
"2310",-0.0109177751115328,-0.0106770913271598,-0.00964897146673926,-0.0170889645734349,0.0110458090817556,0.00578479389715936,-0.0103229748004786,-0.00303019503782953,-0.00462272580999457,-0.0134429144816003
"2311",0.00493963925927043,0.00552767996254167,-0.000885893770173674,0.00620929295989736,-0.00607833387957912,-0.00392588889400591,0.0040639057475218,0.000253183373161159,-0.00829324915751783,0.0151400727276354
"2312",0.000802384995094663,-0.00052356712218915,-0.00443256538921322,0.00154267643704076,-0.00410218208923485,-0.00357447107183906,-0.00256348691674158,0.00177245340906151,0.0160561796946617,-0.00149140393515124
"2313",0.0161371620055348,0.0267155274696498,0.0267141845817738,0.0209488579569388,-0.0101043463336172,-0.0028514266246723,0.0236710481465245,0.0245197536952182,-0.0172016131687243,0.00373407885778065
"2314",-0.0012825000821729,-0.00280611652181595,0.00433645562629081,-0.00603510911617133,0.00314080832612995,0.000738051262141992,-0.00132127093141277,-0.00197394554249386,-0.0128967502588812,-0.00892852630190855
"2315",-0.00162950287649644,-0.00946530326270378,-0.0129532190467452,-0.0142681711065537,0.000939248325212194,-0.000184873036157884,-0.000264570115895979,-0.00296664746625774,0.000763519111813382,-0.00825829985097226
"2316",0.00578735786771944,0.010330511349161,0.00174973435444326,0.0200183742214184,0.00297146951225646,0.00525552777002725,0.0127051307519048,0.0126458230362385,0.0222956682120692,0.0174110485764289
"2317",0.00634390810868357,0.00741314311587216,0.00349333287364639,0.0220411699953849,0.00413211525962698,0.00110059594861189,0.0139831166695923,0.0173849307269649,-0.00381457015721265,0.0111607918898995
"2318",0.00392964928679684,-0.000253674639992152,-0.00348117198112596,0.00531754136345408,0.00209657066191071,0.00174077459412958,-0.00386644619788667,-0.00166700714155887,-0.00274697417997938,-0.000735900819623936
"2319",0.00141894956575239,-0.00482235554949773,0.00436675380370932,0.00205696426162327,-0.0076709690122464,-0.00283522507521872,-0.00646893467155729,-0.00121000178908359,-0.00701171935696865,0.00294554370651778
"2320",-0.000537455815223575,-0.00535580402611435,0.00608701516720078,-0.00234592198952699,-0.000234080092412325,-0.00210927126702043,0.000260295694582968,-0.000726986077475011,0.00294215705230449,0.00734219461659547
"2321",-0.00659939485722982,-0.00820514984818832,-0.0129646446915489,-0.0170488352310828,0.0113248110906745,0.00459528251625785,-0.00704819583593375,-0.0106693606514368,-0.0226300984432167,-0.0211371111512028
"2322",-0.000443025333003222,-0.00723877505686166,-0.00612958604727454,-0.0023923536471846,0.00038587781256072,-0.0010061836870775,0.000796178525149571,-0.00661768236141369,-0.00240115768457971,-0.0059567318472874
"2323",0.000590849280810213,0.00416648672540698,0.0149781045824349,0.00329730512232085,0.0013126502581069,0.00146527437107236,0.00768917297569183,0.0032074336039194,0.00232094898442448,0.00299621356440394
"2324",0.00925009123959186,0.0121887104306468,0.0104165034488115,0.0137435983588492,0.0104847908062939,0.00676738548024858,0.0198655309785067,0.0150027404120372,0.0185249059781287,-0.00224052417919829
"2325",0.00438761660153797,0.0107610392935442,-0.00343631147224333,0.010315488432237,-0.010528950633316,-0.00136284971854517,-0.00154761843471996,0.00823817247724534,-0.0139778037390064,-0.00374246393872524
"2326",-0.00242677252870405,-0.00861853331399198,-0.0163794834997236,-0.000875145206503336,0.00709397287428737,0.00363848737823735,0.00594299117120589,-0.00360495295878094,0.00461145182940137,-0.00150268636214512
"2327",0.00681190440396029,-0.00869325667020604,-0.024539764261697,-0.00291972713170574,0.00260837069509257,-0.000290553751806644,0.000642408074281953,-0.00892416902071635,-0.00603535367252084,-0.0173061642997535
"2328",-0.00323814504493736,0.00128951418532397,0,-0.0120059224915666,0.00061223967851598,0.00118058462278192,-0.00141221723345664,-0.00292052775084028,-0.00667064055417776,-0.0137825107354482
"2329",-0.00998760904486939,-0.0190621861805117,-0.0215633676774732,-0.0195613386255007,0.0109359158094946,0.00399034041669655,-0.00565541717950802,-0.00610147597543842,0.0130004474730874,-0.00232932034986943
"2330",0.0109209633963809,0.0152309967243491,0.0165288532648782,0.012091912332892,-0.00726233753861072,-0.00216792350832062,0.00245600906907795,0.00982267562856243,-0.00611934366413924,0.0108950335716682
"2331",-0.0119657914691471,-0.0168132475420067,-0.00541988570411089,-0.0200119881257546,0.0123450263509142,0.00515973339799403,-0.00541568146678761,-0.00851152215939022,0.0142808189792916,-0.00307932878634831
"2332",0.00269685556473198,0.0176269512506628,0.0290642675560357,0.017372774335672,-0.00632290615001363,-0.00153102548697048,0.00570442367492241,0.0129995616117613,-0.00151758703720095,0.0239382940858939
"2333",-0.00234721154205964,0.0018097883590491,-0.00617808805420639,0.0128819130084703,-0.00128791189422439,-0.000180534427907775,-0.00128905941046908,0.00411651392929557,0.0135100819049228,0.00754137452184356
"2334",0.009312791471068,0.0113546974533281,0.0230906337145482,0.0153802064975663,-0.0069024564740181,-0.00396916035279926,0.00684151213304207,0.00795735388839014,0.000166658336804515,0.02170659899314
"2335",0.0101010132141055,0.0137791221530676,0.0277776602480067,0.0177686914057749,0.00351367778834533,0.000724627639278719,-0.0023077788185254,0.00885179373660772,-0.0106622737860324,0.00512828594201653
"2336",0.0000478978023281673,0.00125846893543202,0.00422300718853785,-0.00486539670820263,-0.00479503750014842,-0.00235324896585054,-0.00642519269325414,-0.00545437576630181,-0.0139765600903401,-0.0080175326796712
"2337",-0.00110563021317744,-0.00175965903549635,-0.00925150592395863,-0.00575218522206178,0.0085652270070935,0.00299352536992714,0.00659628733735262,-0.00238422932218652,0.00691654848504375,-0.00367379462428574
"2338",0.00702669483463714,0.00906576110836199,0.00764005706552329,0.00462827656814868,-0.00432186629551223,-0.000994844093821778,0.0042397866863888,0.00693119354725091,-0.0015264586419006,0.00442479420991582
"2339",0.00315415962627563,0.0197154342883619,0.0151643937050379,0.01526058139409,-0.00312228990159391,-0.00162951138098733,0.0010235945560706,0.00593393419749155,0.0156276883918411,0.0212922283683834
"2340",0.000953046333218577,-0.00244730345711486,0.00580891729824384,-0.00453773727451678,-0.0110006454974397,-0.00507854915522643,-0.0140593062278416,0.00259562843593608,-0.00510119576683066,0.0194104523215852
"2341",-0.00537847841287908,-0.00711478769793683,0,-0.0099714512359006,-0.00594812627359975,-0.00164087665713852,-0.0169822438488338,-0.0112967461331043,0.00378244091970714,-0.0042313265506686
"2342",0,-0.00222385697434735,0.0074258433224399,-0.00604325533661298,-0.00256427834331852,-0.00109511721635203,0.0106815873851811,-0.00071418046237659,-0.0128119161415494,-0.00424916097384553
"2343",-0.00172261744312308,-0.00421010194171156,-0.00655202898889595,-0.00636944368385661,-0.00412893684580296,-0.00109692025040464,0.00626319567027567,0.00905202936801897,0.00288407840261318,-0.000711300967053075
"2344",0.00148577516729387,0.00547123603579913,-0.00412197883332865,0.0107808045966029,-0.00453751437247563,-0.0021045192281387,0.00363093132485437,0.00779037948838956,0.00397525152731326,0.0128112856578488
"2345",0.00205825403916493,0.00469950103966776,-0.000827781369678204,0.00605377193917267,0.00998069703891491,0.00550144062727131,-0.000258481495162721,-0.00163977696562023,0.00286439771350633,0.00913564938547906
"2346",-0.0090756914393465,-0.00516989383495758,-0.0455674466412721,-0.0103152415648027,0.00412359025645714,0.00346525383846297,-0.00232625511911277,-0.00633508790306958,0.0189012095186389,0.00557102644813079
"2347",-0.0053988437047674,-0.00247455633378846,-0.00868069463783261,-0.00434269318500169,0.00255752612540827,-0.000363654838552496,-0.00829020096888622,0.000236199322238173,0.0194575066414584,0.00969530142169384
"2348",0.00794848269571258,0.00744211278874052,0.0183887112393841,-0.0026171650094583,-0.0100682435735281,-0.00290400047182116,0.0133228186937451,0.00873431895633314,-0.00331584305190713,-0.0137173754198485
"2349",-0.00870327043227026,-0.0201917588335341,-0.00945808037617057,-0.028279791297329,0.0125955081546183,0.00593495962752266,-0.00219126598506258,-0.0109990804436522,-0.00227198153638397,-0.015299103572847
"2350",-0.0055781599152025,-0.0130686959677399,-0.00868069463783261,-0.0162017724528839,0.00548566179232712,0.00181522340251727,0.0134349615444784,-0.00567888739166234,-0.00609954461694495,0.000706277775116781
"2351",-0.000195025632255041,-0.00483843422569086,0.00525403475306629,-0.00030482639796614,0.0066850598357111,0.00271811168500924,0.00382416321311996,-0.00023814564976965,-0.00114556092910212,-0.00988003858289233
"2352",0.00365900514419182,0.00307066513994769,0.00522648083623678,0.00152533034763147,-0.00427426688847243,-0.00234932735254201,0.00977788470629637,0.00166631949137575,0.0090931432784469,0.00641481120450282
"2353",0.000826325082086132,-0.00127545529173068,-0.000866609144910213,-0.0127932010388226,0.00314279017435348,0.00190208173782924,0.00804833319882592,0.000712748984843969,-0.0205390323104401,-0.0219545936385844
"2354",0.0124339297654348,0.0102170470806375,0.0251518142722733,0.0191297274525142,0.0000763487659314332,-0.000180979976874829,0.00187118503439998,0.0121112647081438,0.00273519266083389,0.0246197266652655
"2355",-0.00935487410079161,-0.00581545787507831,-0.0186124989147007,-0.00242191794204583,0.0056546493335683,0.00153732541648366,-0.0178060160941886,-0.0114969613128802,0.0094230448977588,0.0233216012391908
"2356",0.000290510990919257,-0.00279743818317868,0.00775853988403696,-0.00273134309840006,-0.0045590776323563,-0.0027084518325452,0.00494388309449434,-0.00617133654177004,-0.00786111182784688,0.0013812676985363
"2357",-0.00871420979213711,-0.0102014412384764,-0.0136868900783947,-0.0179549918508574,0.00969395515480209,0.00380179446972728,-0.00807371890976194,-0.0100312548475927,0.00453941054673446,-0.00137936242976755
"2358",0.00986533813057755,0.0123679347004704,0.0138768205965372,0.0120855200304915,-0.00861796713543961,-0.00360708973331392,0.00788522888743404,0.012304234182426,0.000739495528218725,0.0110497861959944
"2359",-0.0093335925288438,-0.00865362915329904,-0.00684350231313391,-0.00459287131670061,0.00167779537861512,-0.00135735040560414,-0.0151418787349298,-0.00166806088745675,0.00344825935677506,0.00751355819875688
"2360",0.000292929712952583,0.00333749729238608,0.000861315018280573,-0.00984313066340958,-0.0142357507901653,-0.00806600213858699,-0.0139653181040404,-0.00405841109412741,-0.0173457943270676,-0.00745752564579838
"2361",-0.00346495063252183,-0.00614124385532078,-0.00688454425001572,-0.00931962515444762,0.00432456577465157,0.00100502972271088,-0.0107848129900555,-0.0105466991428509,-0.001915029174272,-0.00273227328300718
"2362",0.00631732504892035,0.008238951358021,0.00693226976798655,0.0100345330832161,0.000768842618867893,0.000638952672654014,0.00801271611161236,0.00436045790344197,-0.00133481268036673,0.00410953283883031
"2363",-0.00136256106978472,-0.00306427699481671,-0.0043027998229852,-0.001862638567383,0.00222799059996115,0.000638308470055415,0.000912145573492174,-0.000241269706767855,-0.0028401637527371,-0.00545702180239194
"2364",0.0129621462995744,0.0197234908169068,0.00777856460197102,0.010264173550073,-0.00444594904760454,-0.00164065061073071,0.0119774164486852,0.0125455621143131,-0.0173410400266136,0
"2365",0.00678322273155096,0.0113034865670776,0.006861202536671,0.0120074494669211,-0.00377379679268341,-0.000456683888793163,0.00154377544353679,0.00309714132769479,-0.00272804767106449,0.0116597902841575
"2366",0.000286492601629273,0.00372578985327121,-0.000851777389248687,0.00669301777274689,0.00517901351000227,0.00310614191571679,0.00064260816626649,0,-0.00341939639033861,-0.000677887099525876
"2367",0.00429940049349975,-0.00247455633378846,-0.0025574421030945,-0.000302161869570439,-0.00146110030282121,-0.00191239546050315,0.00436443961878297,-0.00118758405819475,-0.00823467990676474,0.00407050060119052
"2368",-0.0019025443981473,-0.00843477060644759,0.00769222704911066,0.00120914497173041,0.0023873535292751,0.00118623956201369,0.00012768511447625,-0.00784759951033498,0.00380552662673783,-0.00608106773660633
"2369",0.00204930667328429,-0.00125091260201982,-0.000848233218477268,-0.000603809348856621,0.00405740058236681,-0.000338032378011222,0.000639089384653735,0.00143804396560121,-0.00103391351083759,0.0101970756409457
"2370",0.0030436351897638,0.00300616476137194,-0.00848894219078444,0.00815699505868439,0.00720764368147608,0.00310449107247224,0.00536370412844311,-0.000957533817978806,-0.00232882521426903,0.00201895364593252
"2371",-0.00298715754513235,0.00549438081973874,0.00428083357871412,0.0152832779186429,0.0142353271006352,0.00928335475550668,0.00304885223628393,0.0162911614336783,0.0277513534667821,0.00671589392978178
"2372",0.00508842782499141,0.00322901228006756,0.0102301108841361,0.0106257630771114,-0.00743100334555169,-0.00261507305119835,-0.00620557496067964,0.00660097921507052,0.000336482175382402,0.0120079785873621
"2373",0.0015614115706597,0.00693252876816453,0.00675110073940544,0.00905362564034551,0.00242035849388489,0.00144667119024566,0.006117130292147,0.00491805913328647,-0.00084088464246368,0.00988800541244195
"2374",0.00325977510892872,0.00221292091027148,0.00586752742742158,0.00723600182361728,0.00535617924524101,0.00117356064199114,0.00531974703930826,0.0046610226131325,0.0148123379902374,0.0169711811449773
"2375",-0.00136556421526135,-0.0144751519655213,-0.0116667123436496,-0.0114941088173087,0.00645252336844404,0.0015330964739324,0.00151189105520677,-0.0034797268963217,0.00555646034903878,-0.00192551936769392
"2376",-0.00947770285034766,-0.0343538928110562,-0.017706590418109,-0.0252907718399699,0.00484604054526083,0.0035114727893939,-0.00490615991269705,-0.0188545241702737,0.00404122061855672,-0.0122186152959649
"2377",-0.00771157217611829,-0.015210089101762,-0.0180257652605508,-0.0140172981463198,0.00445202423958135,0.00197409185211117,-0.00075874987894009,-0.00972741850252545,0.00739281267279135,0
"2378",-0.00196706829564419,-0.0185863823271325,-0.00437047792040235,-0.00332739140944815,-0.000738912326562313,-0.000268657836696051,-0.00544019915890348,-0.0129370563841105,0.00105999674706458,-0.00651046168649383
"2379",-0.00139375372568873,0.00533458610411208,0.0096575357121107,0.0106222252565686,0.00384420470298674,0.00304566172674159,0.00915913548395597,0.00339806602128201,0.00741225887624641,-0.00524239253493219
"2380",0.00298425008147296,0.00716387433483723,-0.00434776817051308,-0.00360369947819006,0.00485992958107673,0.00107152153710754,0.00504198591712224,-0.000725631330227405,-0.0105110203751617,-0.0171278363614298
"2381",-0.00372415510174384,0.0150156632196461,-0.00174667813171003,0.0027125086425468,-0.00622899003185962,-0.0033896605468785,-0.00150495017695096,0.00383258454009994,0.012828893924552,0.0234584695446547
"2382",0.00644000911454712,0.0254346856002265,0.0227470386524538,0.0177336604622242,-0.0106926305460134,-0.00429657171380982,0.00188432832658547,0.0248055572579324,-0.0059701332626898,0.00916831322138223
"2383",0.00283870414638709,0.0102058203887767,0.00684347940355923,0.00767884428715715,-0.00462124294218746,-0.00224736917046253,0.00411158834686809,0.00783091726152207,-0.0192354761726765,-0.00778717815876662
"2384",-0.00163118826793407,0.00205139537026122,-0.00924826050729399,0.00254016305047422,0.00164739042070039,0.00198212743277537,-0.000503839041888443,-0.00306085714223359,0.000496573998562511,-0.0058862543246091
"2385",0.0130224852533258,0.0307061911943531,0.0224719542385388,0.0241601215488481,-0.0114379725564427,-0.00476602026167472,0.00668083972931899,0.0174775197856381,-0.00653433405236836,0.00789483252926959
"2386",-0.0359091449280415,-0.109483705822347,-0.041419977593303,-0.0607017960977838,0.0268468524805718,0.0138239525775041,-0.0121463438080635,-0.0733520096302124,0.0490383727496597,-0.0202349783501855
"2387",-0.0179097368218786,-0.0231391774433878,-0.00529105252705953,-0.0128637641372736,0.0249668765698479,0.00864425781270195,-0.00190124438439621,-0.0230462026643503,0.00539682539682551,-0.00199870871444952
"2388",0.0180361689679667,0.0322488578113547,0.0150707981251978,0.0294756818776525,0.00208405691223268,-0.000176338111656849,0.0217168282195648,0.0358976233672774,-0.0107357120303128,0.0160213488817786
"2389",0.0170274143236426,0.0221179064701433,0.0131006486853331,0.0253166034108148,-0.00767245260920879,-0.00406538412752677,0.0128032468037771,0.0175741942887906,0.00414934567507186,0.014454602712451
"2390",0.013645362615873,0.0221800393482223,-0.0086208349952257,0.00999407246928352,0.00368498284049279,0.00221854225184548,0.0111682838963645,0.00827049982926975,0.00500639717121421,-0.00582893627845582
"2391",0.0021006683270377,0,-0.00173905372269767,0.0096039923891782,0.013884981364374,0.00264168182176472,-0.000728317622743169,0.000482430122212829,0.0153396298304764,0.0123778149562057
"2392",-0.00719334195837484,-0.0283141997517737,0,-0.021331632949757,0.0125200849119114,0.00548246249289952,0.00765216545751946,-0.0217022242036815,0.00825478519570799,-0.0283139731648793
"2393",0.00599786117963519,-0.00408509899924048,0,-0.0026510535897456,0.00161590421462288,0.000175838353225766,-0.00361603493281459,-0.00147902742305972,0.00587004706982275,0.0039734554960511
"2394",-0.000620001659292324,-0.00519554323595139,0.000870972210665011,-0.00265797223186004,-0.0000698105980287966,-0.00131872134024202,-0.00883146184924688,-0.00271535774487286,-0.00376250491476637,-0.0283641363814513
"2395",0.0148903130464928,0.0156680336541262,0.00696252364129535,0.021616946159615,0.00736572421153592,0.00193682381108506,0.0147685619880022,0.0168318200985744,0.0060120161086783,0.0101833702572474
"2396",0.00352711548024232,0.013531988874429,0.0242005784694876,0.00956517657802114,-0.0087746336601765,-0.00527218873315949,0.00721684904715825,0.0131449388808336,-0.00942392707864148,-0.00403234117737061
"2397",0.00726334840115084,0.0149531247608754,0.00590718166245208,0.0140684309651711,-0.016439435386972,-0.00591893283652367,0.00119401394979546,0.0093704716700127,-0.0165518687900309,0.0188934773809963
"2398",-0.00013954270526273,0.000263106797830481,-0.00167786753442245,-0.00169886693789389,0.0117855648456169,0.00257707557268327,0.00417470025237732,-0.00214225345008801,0.00920176941876893,-0.0125828817108378
"2399",0.00558332368273051,0.0105207224202584,0.00168068750542338,0.0144640663455848,-0.0145431292262506,-0.00416578582375227,-0.00736428475151807,0.00620215308523298,-0.00771512582601408,0.00402422820351811
"2400",-0.00134180518389571,-0.00598662061130439,-0.00335573506884468,-0.00223673022175508,-0.00859617229311238,-0.00382727847991082,0.000837629381511551,-0.0111428405715059,-0.00384831534048036,-0.00267204288248979
"2401",0.00268729045881577,0.00235677197765916,0.00252532019097984,0.00896612671306074,-0.000939367600925167,-0.000268345986797702,0.00251081213674675,0.00311687315548026,0.00157682912572787,-0.00468862042717499
"2402",-0.00101669962209661,-0.00940454906721933,-0.006717105044455,-0.0102749197932618,0.005640808506018,0.0026813821327849,0.00453191168432654,-0.00286793353732362,0.00133814545546174,-0.00605644537272443
"2403",0.00416300828359684,0.00870269836215631,0.00845313962173666,0.00505078031578177,-0.00546589419620702,-0.00204970558826578,-0.000237531979495387,0.0105464478463173,-0.0143070514449103,-0.00677045791683872
"2404",-0.003777119687563,-0.00235284467865982,-0.00754400793799903,-0.00307119943309142,0.00202497288489378,0.00223265598339761,0.00142504599625037,-0.00189743349768268,0.0152325067009531,-0.00545330161916657
"2405",0.00448520723456691,0.00183427731537855,0.00168920442888099,0.00728079145209581,0.00173236846254099,-0.000802295843780776,0.00830068375236315,-0.0007128864521736,-0.00746272566859252,-0.0020562452815841
"2406",-0.0027159248181593,-0.00026159272880999,-0.00337271165829134,-0.0100081329403624,-0.000720344560005026,-0.000802652174884178,-0.000940908882927527,0.00356721664112158,-0.0069647567386586,-0.0109890024443174
"2407",0.000461550137214273,0.0034015089598014,0.000845986373307017,0.00786289343782021,0.00158619709801999,0.000625032992947361,-0.00459069544135193,0.00545005115063724,0.00422410931518202,-0.00416660978580086
"2408",-0.00106113235142158,0.00651872272929421,0.00169063241664791,0.00334350013311635,0.0124530328714343,0.00428172779210012,-0.00709565648130994,-0.000235688618740904,0.0161111031746033,-0.00976298245846985
"2409",0.00115471890524721,-0.000518027998477111,0,0.000277573548180587,-0.00184867989223181,0.000532742969874711,0.00738436351381533,0.00495050808751873,-0.00288990863774041,-0.00281693550467965
"2410",0.00161452369946491,0.00959049530291134,0.0177215898345422,0.00527502341301633,0.00833439322257923,0.00381786541182727,0.0096951624159185,0.00680272473505661,0.010339902543008,0.00847467913859545
"2411",-0.000828898212204443,-0.0107833181597822,0.00331669126886069,-0.00193312148470437,-0.0108423374014669,-0.00347217068342021,0.00351282544434905,-0.00582485766780061,0.00186079242861803,-0.0175070513551416
"2412",-0.00640744112200575,-0.00259518860705998,-0.0123966526536556,-0.00719428260298793,-0.0103025917291484,-0.00239931895204082,-0.015169151644571,-0.000937362690721644,0.00812570029309945,-0.0014254239409307
"2413",0.00292258755625752,-0.00416341496780404,-0.00502094348233828,0.00334455287821367,0.000577964701123035,0.00053466320328921,-0.00426531179581102,-0.00821022199426058,-0.00475942259125139,0.0164167665089441
"2414",0.00106407891492188,0.00418082146245857,0.0142977688808279,0.00555548274859063,0.00751405483692924,0.00240393822522367,-0.00238013671474857,0.00709550371073986,0.00169688399677059,0.0042135701416901
"2415",0.00817887603849865,0.00338280686464532,0.00331669126886069,0.0116020827033498,-0.0103974725758902,-0.00621761110178665,0.00131192197298979,0.00234858359270018,-0.0178639569517192,0.00419567454347969
"2416",-0.000596016037349045,0.00103724475521405,0.00413229075220345,0.00710010252797888,0.00188369774883523,-0.000536431282646688,0.000953108150856474,0.00234305092602693,-0.000862414719033699,0.00557102644813079
"2417",0.000596371484318015,0.00958532766417997,0.00905351371033092,0.00677866801818694,0.00983649812740506,0.00357704229205646,0.00368916030302913,-0.00233757387140299,0.00408032793345359,-0.00277004539170966
"2418",-0.00247499116050065,0.00384923998258291,0.00326258532122714,0.000269317577300754,0.00386755039592845,0.00267313094467214,-0.00130414431516357,0.00421748571767844,0.00468895752335863,-0.0118056088131202
"2419",0.00464070987308718,0.00792437671770929,0.00731716084817857,0.0129240551367171,-0.00891808170317299,-0.00479855197200874,-0.00949780782766774,0.000233353647363765,-0.0069228376932613,0.0154603742383221
"2420",-0.00086895076213056,-0.000760838736615588,-0.00484272265898678,-0.00372139381394476,0.00842235347063935,0.00357163292460005,0.0027568464675729,-0.00186603828097043,-0.00211479599145925,0.00761242387006322
"2421",0.00288380411465305,0.0020303457663291,0.00567719679079715,0.0104055619487864,-0.00942299494122023,-0.00293634275962529,-0.000717261382575662,0.00397284848346757,0.00345364201799625,0.0164835036664763
"2422",-0.00515762950186605,0.000506592783606541,-0.00887098386552854,-0.00448899164311867,-0.00266637681508997,-0.00169571463800677,-0.0117224129405556,-0.00256070802745056,0.00492807430938913,0.00810813667656118
"2423",0.00188109730754826,-0.00151889743291322,0.00813683525078801,-0.00636621200819987,0.00599723414907949,0.00160935143199725,0.00290474884090952,-0.000233171112013264,0.000233509767000095,0.0040214617765566
"2424",0.00224380897685394,0.00760676515409209,-0.00484272265898678,0.00934333827268596,0.00158045297666698,0.00178510970498502,-0.0028963357131041,0.00373454173576127,0.00474708949416347,0.0126835420999869
"2425",-0.00146220783364515,-0.00830413183901324,-0.00243306894558803,-0.00555404020045069,-0.00523490966555562,-0.00338583120634672,-0.00726236591588714,-0.00697646006431718,-0.00882968004934037,-0.00329593395865624
"2426",-0.0000456505812552743,0,0.00569097868233404,-0.0132977285756044,0.00843492121708844,0.00223504544769448,0.00512090501041995,-0.00210787380776523,-0.00148473859900955,-0.00925926871340432
"2427",0.0020133741106354,0.00456729280295476,0.000808522205114404,-0.00404308823159705,0.00107161764190233,-0.0000891978465831222,0.00218340767433123,0.00657122504796659,-0.000156495540432733,0.00400528569093561
"2428",-0.00511474875317075,-0.00303097200975255,-0.000807869025068797,0.0027062069080499,-0.00235592131000339,-0.000356669873750159,-0.00484144467915837,-0.00373072145830999,-0.0111146366450433,-0.0119681274213354
"2429",-0.000688656519483799,-0.00430711468522693,-0.00485031695385063,0.000809843647337827,-0.00379440392804586,-0.00160632531061,0.00364859365696169,0.000468305601582175,-0.000870611077112948,0.00403776877017403
"2430",-0.00188334907005894,-0.00534354409997706,-0.00731113005757034,-0.0086302502180553,-0.00581977865725114,-0.00384369919432659,-0.00933103968232596,-0.0112279558466417,-0.00142596843636289,-0.00335122964418233
"2431",0.00492442278476779,0.0046046820101846,0.00327333007381103,0.00761700081702932,0.0133710390645683,0.00412763136837135,0.00941892807394895,0.000709652076160472,0.00198333989726285,-0.00403491472006745
"2432",-0.00164868119691464,-0.0015278773751648,0,-0.00269963206214296,-0.00385162483043011,-0.0000893572535060061,-0.00169647900710401,-0.00520084491595263,-0.0100554550263946,-0.00945308182100768
"2433",-0.00284419919178325,-0.00178515773026822,0.00163133600801246,-0.0110990785711613,0.00143149100641282,-0.00116194972523653,0.00194224191687731,-0.00166363302491657,-0.00199952013116467,-0.0190865205881448
"2434",0.0000461944719336582,0.00562087054085847,0.0073288394992892,0.00766495756642405,0.00110351271160414,0.00156824854673832,-0.00169619133811594,0.00928360195463407,0.00408720952145547,-0.0111189659261556
"2435",0.00450806995996977,0.0149899206838155,0.00727566875950036,0.0162998820965412,-0.00815671655373507,-0.00259438292468928,0.00800968313333894,0.00117909716052234,0.0102162901251792,0.0112439874393682
"2436",0.00302234972146875,0.0055066019856127,0.00561796470864251,0.0213846385064682,0.00728621434619536,0.00466380644093367,0.00710326533669137,0.0148411192570523,0.0169076953464486,0.00694917489634173
"2437",-0.0000914682029690139,-0.000248959210288557,0.00478861486759019,-0.00314060607949462,-0.000716266212181904,0.000535448874200206,0.00573835790535737,-0.00580298803461199,-0.00341856092044179,0.00897172432975935
"2438",-0.00228280508871437,0,-0.00476579331884763,-0.00262512764873257,-0.0125413771872306,-0.00490717659872286,-0.0114110320028225,-0.00256859867298997,-0.00530137973645028,0.0177838964431223
"2439",-0.0239348802104161,-0.0209161378150358,-0.0159616254252044,-0.0336934662592854,-0.0164740776300769,-0.00475202201949887,-0.0397979219810228,-0.0255147462354648,-0.00658355691146817,-0.0154570542315235
"2440",0.0143473036928281,0.00890115298939409,0.00811035193900511,0.00681038613873675,0.000516318649557368,0.000900963377244102,0.0121462160880474,0.00480432527422026,-0.001262358974359,0
"2441",-0.0143754734088218,-0.019914088996399,-0.0176991460696774,-0.0251624115476015,-0.0113578448760638,-0.00369056099522624,-0.0243723232515276,-0.0207987795299202,-0.00663556384028952,-0.0129693172763443
"2442",-0.000375378152123296,-0.000514495334514309,-0.0065520439634662,0.00305311929690544,0.0014920917890644,0.00225841640026947,0.00304346196532657,-0.00170875134537429,0.00341948310139162,-0.00760708883651384
"2443",0.00999310386074304,0.00797728238558837,0.00494652442731858,0.0171553061071559,-0.00432075262990872,0.000270485555225131,0.00455121933097002,0.00611378563747511,-0.00641937708036144,0.00487798195622902
"2444",-0.00386553706571002,-0.0178708184435823,-0.00820358433658464,-0.00680067968146369,0.00807979930586877,0.00108147562729033,-0.00100686488020207,-0.0110592129160868,-0.00247272068741999,0.00138694364428016
"2445",0.000187459043390126,0.00779833701170252,0.00330854954204374,0.00794292848013511,-0.00326507413086474,-0.00170998597991712,0.00944821346598923,0.00793491155760218,0.002079018104574,-0.00069244007257252
"2446",0.0000468173120782289,0.00206333820365767,0.0140148787192746,0.000543494790867349,0.00349930368703366,0.00153282305982239,-0.00162203831377083,0.00442772368007427,0.000957564634535668,0.00346495601403118
"2447",0.0112454818033434,0.0128701099524231,0.0292683193444581,0.0279741737341372,0.00808731941672791,0.00162053983407962,0.0114996166818049,0.00857214400104644,0.0145886078668909,0.0124309117376125
"2448",0.00630142661406041,0.0116901260993136,0.0126381345563149,0.00713313508244195,0.00794859900413147,0.00296617162742607,0.0194021761789969,0.011413245159847,0.00235721699592717,0.00545709200812983
"2449",-0.00547927591569286,-0.00753595493055881,-0.0140404821098483,-0.0128540097729919,-0.000949019022029485,0.0004481400701557,0.00254560919782532,-0.00408135541065358,0.000627122364192267,-0.0115332945108013
"2450",-0.00810199169684189,-0.0111363548469304,-0.0087026311513686,-0.0146159364462848,0.00635874691749416,0.00286676173972644,0.00117065889680767,0,-0.000783384241545115,0.00686346568920571
"2451",0.00620783614560771,0.000767736603415781,0.0111732650376719,0.0142933693063589,0.00733511388635666,0.00169692610859551,-0.00779521685823192,0.0077145865414614,-0.0072912581585749,-0.00954336553088786
"2452",0.00496355976176166,0.0112533555499574,-0.00157854623374787,0.00904016321940171,-0.00216289058860364,-0.000445758696838938,0.00552413118532735,0.00334910691235013,-0.00315907432098228,0.0233998982825621
"2453",-0.00904740615102051,-0.0144160519769228,-0.00711470992276098,-0.017391345103953,0.00252883408329807,0.000624424708573601,-0.0107435916991464,-0.0164521673951005,-0.00118840911750584,0.00605251050862865
"2454",0.00754609942950668,0.0105210771718134,-0.00159220199293086,0.00429076648435722,-0.00893700765032179,-0.00249636018615274,-0.00481289659576856,0.0111517012790889,-0.00341081145395405,0.00334226902923129
"2455",-0.00240389281014008,-0.0015235257188092,-0.00318982132203227,0.00694251052310624,-0.00330014993025884,-0.00232708493169098,-0.0181052328458281,-0.00455530885919142,-0.00254695162804008,0.0086608425336514
"2456",-0.0050979443985556,0.00152585039112307,-0.00559998670126716,-0.0111376219313902,-0.0116954567206429,-0.00457529118997657,-0.014397498299806,-0.0139690956646316,-0.0347111315033514,-0.0026419718257199
"2457",0.00442534625574842,0.00253925608903294,0.00643607838030191,0.0144810678501628,-0.00465928608741228,-0.00225292268153821,-0.0193491382264798,-0.0134344432662343,-0.0015706538681437,0.00596018324407677
"2458",0.000695641893207588,-0.00607894622013694,-0.00479626978176939,0.000793117151379086,-0.00557270946618971,-0.00207756024925687,0.00169870083247559,-0.0118842176087091,-0.00927301713258011,0.0019750244006882
"2459",-0.00342927135478843,-0.00764519932650454,0,-0.00449040595762129,0.000672432616404262,0.00144839592621682,-0.00143502058280365,-0.00876952752210725,0.000668510758197849,-0.00262808499404299
"2460",0.0052081838935838,0.00231137933535108,0.00321294457740495,0.0108783322451635,-0.00589849231673556,-0.00262145647004364,0.00587847073529746,0,0.00350764996672215,0.011198928205062
"2461",-0.012629704839679,-0.0148605701018741,-0.00880706088130723,-0.0230972152953798,-0.00225394595062334,-0.000271703066453188,-0.00999998774074917,-0.0171891492920493,-0.00507657273380246,-0.00586324608441957
"2462",0.00131207909142672,-0.00286076982234174,-0.00161552341398208,-0.00188057710350076,0.000978885198557045,0,0.0135118879352345,-0.0015432495375397,0.00158925131938314,-0.00720842462624149
"2463",-0.00327540128398673,-0.00443403052218161,-0.0016181160547396,-0.0088830156201829,0.0037603821598331,0.00208468156315056,0.00556565964219335,0.0108193790281232,0.00242192253920037,0.00660070625287879
"2464",0.000516347340260737,0.00104795810427083,0,0.00162962815027989,-0.0140116646337585,-0.00307545566956435,-0.00334668885458977,-0.00280334423155726,-0.00558192123287449,0.000655728765314612
"2465",-0.00347215280078161,-0.00366421516198645,0.000810401598727362,-0.00108457276699547,0.00638370713431158,0.00217776599438069,0.00129142210795297,-0.00536676726098939,0.00268095674697588,0.00131066557908799
"2466",0.00626228441146459,0.0123461006777812,0.00566785189063124,0.0176437963425582,0.00324639510955271,0.00199172277253767,0.00683601956988245,0.0125898198868435,0.00618313836898388,0.00196339129656375
"2467",0.00266701283303261,0.00155661728325573,0.00322064133799782,0.00613488076135904,0.000828220422389947,0.000451732353058398,0.00422773615814509,0.00558224912985317,0.00572997019980015,0.00653165629159558
"2468",-0.00186656016735876,0.00025917074424564,0.00882833079239864,-0.00291606920989806,0.00105303889215791,-0.000903134180424647,-0.00382724993178063,0.00252368134458325,-0.00305509864540421,-0.00908501892228064
"2469",0.000467378273863117,-0.00259012418709259,0,-0.000265995717653622,0.00150273428020498,0.0010849150224479,-0.00128060817814868,-0.00226544352566371,0.000745436487418205,0.00392921932243606
"2470",0.00425296806677955,-0.00129836804460626,0.00159110425844444,0.00425527545179527,-0.00435093892250837,-0.00135464020918974,0.0026927989867529,0.00227058741321851,-0.00223457746859923,0.000652373967855002
"2471",-0.00335070722214059,-0.00260002618303401,0.000794246122462594,0.00105952662299025,0.00263700428008473,-0.000180645393306089,-0.0019182171886768,0.00125822074561532,0.0075481338345742,-0.00456323801298775
"2472",-0.00200762639419994,-0.00547437144167284,-0.00158737921437313,-0.0105820149845479,-0.00676313681821894,-0.00217068482943095,-0.0116591620404904,-0.0103064568884379,-0.00559809001730394,-0.00654883367309145
"2473",-0.00266686755471557,0.00183475815514944,0.0015899029933375,-0.00855614753053668,-0.0108939502800435,-0.00344424463007864,-0.0229453376677956,-0.0111760628425183,0.00182135109014525,0.0059327489710721
"2474",-0.00295537372932297,-0.00130821954003113,0.00158740030322813,-0.00404550291354611,-0.00221816703116351,0.000181921013402198,0.0019901234554649,-0.00616493984473665,0.00471035443830492,-0.00655305811402018
"2475",0.0000470840944069018,-0.00104784282369175,0.0007923580068534,0.0056864747327996,0.00613286287887438,0.000818685642922423,0.0148307473799931,0.00749554963937826,0.00296101327585108,-0.0131925678921104
"2476",-0.00724542458348565,-0.00445856586976356,-0.00395896894499981,-0.00807743955302287,0.0000759207715539389,0.0000362426914586322,-0.0220513984972407,-0.00384825784296094,0.00647860412533041,0.00467914912177814
"2477",-0.00601860770774543,-0.00711277778487773,-0.00635918952566294,-0.0119434304052429,0.00435126085665472,0.00300221316740479,-0.012808413622535,0.000772715575718674,0.00741461727170334,-0.011976089318696
"2478",-0.00457713088434242,-0.0021224920765549,0.00239989408630681,-0.00274745485220673,-0.00767637043196079,-0.000634863678568132,-0.0058116351899693,0.00257329802696771,0.0053381106869792,-0.00336702670285538
"2479",-0.001101473318733,-0.0090403046697155,-0.0119711448455531,-0.0101928334653643,0.00896080949714029,0.00308595986638127,0.00530176738259192,-0.00770027329177136,0.000724022508671984,-0.00675673420271494
"2480",0.0220566527172301,0.0160987306482849,0.007067796886286,0.0361814463486601,-0.00850192416143059,-0.0041623550035409,0.0163624992677296,0.00931189643035979,-0.0180078544738954,0.00408164694177549
"2481",0.00450398651706729,0.00316886716477427,-0.00120309639231997,0.00644643535599121,-0.0040570753776773,-0.00354379291851759,0.00612030030827726,0.00256274673815016,-0.0041752189246792,-0.00135499503103398
"2482",0.0106021399718841,0.00500134286684317,-0.00843211777843456,-0.0325594726249419,-0.0424324942601815,-0.0152288311235224,-0.0185134777213687,-0.00434537210648578,-0.000657686621651554,0.00474898719275374
"2483",0.00249565329653212,-0.00366674856166804,0.000809995506815708,-0.0284137164936527,-0.0147705107421705,-0.00601918046070438,-0.0181893718844762,-0.0269578417287293,-0.0148897501627139,-0.00810266141648341
"2484",-0.00230504442292723,-0.00972678224885215,0.00141610299859818,-0.0190233215188182,-0.00562222337313001,-0.00204960227281903,0.0053520926194206,-0.00765169066578553,-0.0221294530271399,-0.0190606052729353
"2485",0.000785434958517905,-0.0082292863702822,0.00121219656033267,-0.0072358120129743,-0.00598175317858618,-0.00578794416446193,0.0169259851081727,-0.0124964736114712,-0.0084542870786386,-0.00208185917709702
"2486",0.00780291567272506,0.00588867460786324,0.0016142194400377,0.0201166437499278,0.00494590637662129,0,-0.00362417821704242,0.00700049122509072,0.00869866498407834,0.0222531114282418
"2487",-0.00187850331989214,-0.0119745195932006,-0.00483485380511139,-0.00828807021708278,0.00902333808099365,0.000938912537956194,-0.00215560530955816,-0.0131017260714167,-0.00298843913110214,-0.0122448708106266
"2488",0.00514075906773126,0.00457852786953694,0.0149798054214234,0.00144098150397109,-0.014714252902833,-0.0044090606365198,-0.00823552469114452,0.0149008684632426,-0.00513829763993223,0.00206601655464245
"2489",-0.00223770473503282,-0.0109920081903816,-0.0149582825618577,-0.0046045807107481,-0.00288789733764239,-0.00442828410808216,0.00299494169709269,-0.00854203962192956,-0.00878020158010162,0.0082475228783081
"2490",0.00755164522720664,0.00975890952754099,0.00809885754243034,0.00982963644135126,0.0024825008192646,0.000851739109619443,0.000135910241953807,0.00215384090955228,0.00373425959645224,0.0279482321863713
"2491",0.00195331508040342,0.0010737223278694,0.0024100802617204,0.0151731823314931,-0.000330158317275342,0.000945965986584252,0.0170984058039132,0.00537343536420498,-0.000346089282815432,-0.00132631000327676
"2492",0.000543994942349801,-0.0072404863779717,0,-0.0107161969996484,-0.00388086346216043,-0.00359040223148532,-0.00547008771526969,-0.00213785944670508,-0.0198199842494375,0.00398407763104802
"2493",0.00371543929323814,0.00810378146257595,-0.00841513851374687,0.0048458880349993,0.001492213954287,-0.000853192439144279,0.00509784115262457,0.001339024801011,-0.00565120529801322,-0.00727510080633487
"2494",-0.00469492454281717,-0.0112542053455486,0.00868852025258904,0.00397172123160461,0.00736634936997849,0.00455522677148013,0.00347053050476265,0.0074885788990231,0.0105674628312986,0.00333106690960094
"2495",0.00195039153523946,0.00840124719349267,0.00100168627622743,0.00141267212497809,0.00419023670349472,0.0010388149381757,0.00824657393124362,0.00398201761282935,-0.00465734609866397,-0.0199203198141998
"2496",-0.00239917696510583,-0.00080611308483225,-0.00160095386365633,0.00169311506731318,-0.0162005012916275,-0.00669986129785782,-0.0125327932107059,0.00026453916395841,-0.0134192375762137,0.0304878065787826
"2497",-0.0036754976740323,-0.00134504952539805,-0.00841844810814474,-0.0118308563777816,-0.0105585078141616,-0.00381508788866347,-0.0157647266858393,-0.0129528032920327,-0.00187918568232659,0.0184088928598929
"2498",0.000500920701579144,0.0029627981907856,0.00303211430700312,0.00114013074727692,0.00732760136413857,0.0044884309555715,0.0105873487658346,0.00723080133169107,0.00537921816945297,0.00710139187360448
"2499",0.00600878040723218,0.0158430586950693,-0.00120909367134381,0.00825742224405102,-0.00108671153245488,-0.000380359632394023,0.00792517565032202,0.00452006801584104,-0.00535043700151983,0.00512820106818124
"2500",0.00316742995069585,0.00978054477025436,0.00443891044348366,0.00536589399916698,-0.000753479023549719,0.000380504360892875,0.00639629172143596,0.00608797828815155,-0.00098620225043744,-0.00446429040277008
"2501",0.0130807670587083,0.0141361795103181,0.0148655216547371,0.016853740206477,0.00854409109492993,0.00332769222092888,0.0194650862297432,0.0142067875567915,0.0035897155164677,-0.0076874068323729
"2502",0.00244865889846535,-0.0043882478091134,0.0114805365683655,0.00441984388323546,-0.0117941311848104,-0.00379052551968118,0.00506545042220208,-0.000778197414300519,-0.00232497536752252,0.00193683988393856
"2503",0.00604051998695798,0.00518530702376729,0.00293545770326764,-0.00522557698395609,-0.0124389773692943,-0.00513622539009284,-0.00077526409271178,0.000778803477152756,-0.0104866720444563,0.0051545684159735
"2504",-0.00114787632022562,-0.0015476100557229,-0.00975616473538754,-0.00663526532740355,0.00187231940383703,0.000191257703630932,0.00620813106502416,-0.00544738190010352,0.00380432964122579,0.00641030081676885
"2505",0.00667399911989852,0.011624881770014,0.0118225998887822,0.0111328850754264,0.00356767598598839,0.000573183374487529,0,0.00808548328691128,-0.00333877458942422,0.00254773579355727
"2506",-0.00825416211693453,-0.0145556632179705,-0.0153844972427879,-0.0297276510480933,-0.0111732714616283,-0.00831174647483435,-0.0185090361206495,-0.0165588839622253,-0.0146672253870682,-0.00952992615734338
"2507",0.00411715741253449,-0.000259009857141002,0,0.00170233326853575,0.00505078482902843,-0.00279356680907328,-0.00746477787108146,-0.0144701699046251,-0.013691132708056,-0.00128285619031576
"2508",-0.00195576840565537,0.0031103207068246,-0.0087026311513686,-0.00453133898924696,-0.00229948818787806,0.00125603767999505,0.0133265380589018,0.000739597435251538,0.00661456145386863,0.00449589628991709
"2509",0.00217735422727694,-0.0036174797307349,0.00857937101521333,-0.00682793280413396,0.0107562142364808,0.00463111518797144,0.0110678208195145,0,0.00499762133278225,-0.00575452855061109
"2510",0.00385747447642881,0.00363061340112347,0.000989223359052493,0.0034373593216559,-0.00498316299395207,-0.00211265459446219,0.00180272627380518,0.00653396135813189,-0.00736711510699384,0.00450167871434171
"2511",-0.00278256250420483,0.00155038094225879,-0.00533814874620586,-0.00415763230108601,0.00441406976685865,0.00163597747016264,-0.0123055321443966,0.000282194720494067,0.000556610069982311,-0.00576196249489347
"2512",-0.00172742037483742,-0.00179365080311122,-0.0016080689218011,-0.0118875843928827,-0.00178802321120775,-0.00043305754074352,-0.00184768760787213,-0.0039503117303602,-0.00241077426816461,-0.00128774623731354
"2513",0.0014643299499002,0.00286456900604581,0.00181188029469825,0.00586845449117535,0.00203709364702309,0.000962797835891926,0.00264440214459971,0.00481581439775924,0.00316018229055426,0.00193420953618118
"2514",0.00248087389180629,0.00129848645526942,-0.00622978850052258,0.00437589709957065,-0.00321890149657622,-0.00144315135628548,0.0011868030170199,0.00535661975532209,0.00583709811915112,0.015444003425422
"2515",-0.00826447695969956,-0.00622414269811666,-0.00141551688143693,0.00755131276155319,0.00730861583526488,0.00366079178270806,-0.00592699552347153,-0.00701062537397512,0.00276347646948194,0.000633704922959666
"2516",-0.000222761089029189,0.00704599457521748,-0.0101255988208752,0.0164313849511095,0.00354343007647717,0.00307130148832102,0.00993756638566001,0.0104490047959822,0.0131361380384334,0.00126673755373652
"2517",-0.00365495263330695,0.00570092973534786,-0.000409140361173121,-0.00709021535865395,0.00151314819704407,0.0029661072869942,0.00944632243221588,0.00838471377715866,-0.00616556345846808,0.0018974420434541
"2518",0.007650020598444,0.00231906770749335,0.0081866295744395,0.0119965726440947,0.00428125534063151,-0.000476862884361218,0.00402906015305682,0.00083120145340887,0.00784599938102359,-0.0119949157764663
"2519",0.00594916160736991,0.00874022816271225,0.0200973794707395,0.00762080112462349,0.00384493229557648,0.00114527554619803,0.0137218083916817,0.0105237236769467,0.00353037020430547,0.00766769250680732
"2520",-0.000794581021897778,0.0086647767071828,0.00577122146174802,0.0109242761796342,0.0156533337808724,0.00648327056763076,0.00344788039494692,0.0150725665131373,0.0155150729251752,0.00507298460463712
"2521",0.00357784551588325,-0.00429517165032223,-0.00158307836347038,-0.00415628647354194,-0.00918176717594488,-0.00454703278304014,-0.00216346967824688,-0.000270056298044663,-0.00737255272033122,-0.00126187729913718
"2522",-0.00330079961172036,-0.00380622194144142,0.000991083888692623,-0.000834726657825358,0.00802561057834783,0.00380631956926969,-0.00663195278870399,-0.00189023459951354,0.00823264429530202,-0.0151611396094232
"2523",0,0,-0.00376170351730831,0.00584784861520915,-0.000656513050228402,-0.000473844237934284,-0.00937198419278085,-0.000541409532573978,0.00426026456483997,-0.00448993064839287
"2524",0.00282597534324291,0.00534901484814365,0.00655814060505455,0.0119048329426903,0.0033675958017485,0.00113815984612975,-0.00427694670101686,-0.00243606321717282,0.00309322133286405,0.0109535241994081
"2525",-0.00250985117916158,0.00177349993215992,-0.00157941201118128,0.00437761535614389,-0.00221017383147704,0.000568286430022935,0.00455558999121752,-0.00407060808676607,0.0036123700440529,0.0146590152638848
"2526",0.00229549987367972,0.00379359743935348,0.00632768355008784,-0.000817218078311588,-0.00475840690151175,-0.00217743474919396,-0.00103645466739954,-0.00108994290928566,0.00263361416438879,-0.00188439640516536
"2527",-0.00352343118168275,-0.000755846587652598,-0.0112006175049303,-0.000545335604600461,0.0104689824120285,0.00502885954790599,0.00674452008372062,0.000272726636850518,0.0143595045474083,-0.000629382790976241
"2528",0.00220989652564096,-0.00378211914845306,-0.000198642955844042,-0.00545551257239241,-0.0128078352674155,-0.00708100285662949,0.00167456636559504,0.00054536900380886,-0.00845917148828956,-0.008816065726727
"2529",-0.00370452581306357,-0.00253099446464655,-0.00278286955724194,-0.00301697350156638,-0.00685907056022228,-0.00380334280223549,-0.0104179297471921,-0.00981180660684666,-0.000870601526840709,-0.00317664205244783
"2530",0.00367404686467343,0.00532846138402343,0.00637842796997545,0.0019256483845167,-0.00199705635868608,0.000477090391061141,0.00636853766724865,0.00385353778675568,0.00243971427480294,0.0114722499988849
"2531",-0.00260223841753804,0.00328137031188236,0.000594088797734704,0.0148270569749624,0.0100050735392725,0.00524713015227452,0.00761981474438378,0.00795163754755657,0.00643196854153927,0
"2532",0.00641179089666477,0.00201254826811592,0.00257336232983607,0.0062229211077367,-0.0068517820315771,-0.00379590137568697,0.00230709312601252,0.00108826044907162,-0.00449092318429123,0.00252050941723025
"2533",0.00865558028112834,0.0120511733746524,0.0104639001615463,0.0110244592132693,-0.0125505591458194,-0.00495385474871235,-0.00537101525251682,0.000543378159087782,-0.00824149409841668,-0.00628526933019513
"2534",-0.00104545533723555,-0.00620192319802526,0.00136766917038544,-0.00425536829860129,0.00336684145941901,0.00134023971657027,-0.00102823170392008,-0.00461713671283204,-0.009272200839748,0.00442745156679414
"2535",-0.00156975033869566,-0.000499243626010948,-0.00819507373889461,0.000801398748848881,0.00360733485372533,0.00124318790772882,-0.00939511359502099,-0.00136419890175388,0.00203069041090065,-0.00818635137568224
"2536",-0.0062017618166641,-0.00874131828248248,-0.00275431775039814,-0.00533757885371866,-0.00300929361784785,-0.00028668217857919,-0.00688565287171927,-0.00109285644339918,0.00422947403699836,-0.00571427301828686
"2537",-0.0000877993154834167,0.00377917792158833,-0.00236716587615005,0.00187834439384749,0.00695934566743506,0.00343862536987771,0.00784902386147346,0.0095732547204328,0.0138633147857918,0.00574711359443247
"2538",0.000395524708310502,0.00326325038439301,0.00533898429387358,0.000535351875829315,-0.0061833154779849,-0.00191631328294095,-0.0118119426764557,0.00189647610235855,-0.00302904362538192,0.0107936340731034
"2539",0.00065896891815842,-0.00100095402576972,-0.000393367056473082,0.00428281959216603,-0.000419976947245493,0.00038211637185781,0.0111651502232666,-0.002433683553139,0.00555554701967576,0
"2540",0.00689290110201579,0.0040070894933697,0.00452573907890552,0.00612992666580281,-0.000419727420801541,0.000763798451137943,0.0067549332040937,0.00542167856521436,0.00250346175771621,-0.000628132135055082
"2541",-0.00178764469820758,-0.00947872216163737,-0.0015670985090328,-0.00238411216811607,0.0060501308760208,0.00477054406004096,-0.00335486231604287,-0.00188755876837099,0.0135193321325926,-0.00628526933019513
"2542",0.0000437436776030697,-0.00125902747056506,-0.000588638418962173,-0.00504507797170339,0.00735052968085914,0.00180445540706664,-0.00142402895009486,0.00216091566287524,-0.00203906547253352,-0.00442764686394759
"2543",0.00131026949684188,0.00252153205859806,0.00294467809241827,0.00613822140535336,0.0135988425591058,0.00407578533527553,0.00726040268818973,0.00539079969336309,0.00621490725536278,0.00381195738522355
"2544",0.00593250726469363,0.00402391944384473,-0.00137007854487714,0.0045093712544626,-0.0115347369233129,-0.00594740700346286,0.0030892662547588,0.00428948415372377,-0.00761486576504167,0.0050632218761828
"2545",0.00394629345688013,0,0.00705605879750415,0.00924212936540303,-0.000579310110802256,-0.000664665434889966,0.00769905312498387,0.00106786174313389,0.00264299597030426,0.0107053384040592
"2546",0.00544256734895843,0.0045089784226362,0.0038926346481678,0.00313972526534179,-0.00314709850871886,-0.00152064192105461,0.00331097309290329,-0.0029331721212047,-0.00680267868712037,-0.0112149924655612
"2547",0.00399540682278055,0.000748336411536821,-0.00717354722988917,0.00104333670624057,-0.00722688105937264,-0.00361667757083417,-0.00558448023272418,0.000267591595367378,0.00111298798511172,0.00126028713508397
"2548",0.00522024283855904,0.00274107749348462,-0.000976179084352213,0.00807695702322619,-0.00460195705963218,-0.001910530990473,-0.000893535459356221,0.0018717237922099,0.00444707944924305,0.00125863603933829
"2549",-0.000851142336114052,0.00472165339998631,0.0011726581030711,-0.00361836771855262,0.0054639576725366,0.00401960135144397,0.0047266429097661,0.000800272248985934,0.00536402738264852,-0.00628526933019513
"2550",0.0015760881655158,-0.00321562893528105,-0.00058560126906182,-0.00415050131909678,0.00593565194780776,0.0026692461687472,0.00165296063906339,-0.00106672263084584,-0.0033875507556308,-0.00189763734060744
"2551",0.00595519655185961,0.00124089317216436,0.00840010990280105,0.0109404604500907,-0.00174529743412699,-0.000475559745626741,0.012566668894455,-0.00240240501694389,0.000594833446634802,-0.00126734462309919
"2552",-0.000888038539359925,0,0.00116237104316563,0.0030918835432161,0.00166514416760655,0.0016168539133028,-0.00250736788777783,0.00240819046580065,0.00135884501061567,-0.00507620312805912
"2553",0.000677267023284189,0.00272602417953638,-0.000967606015941369,0.000256826045995195,0.00299239710724675,0.00265894565994418,0.0042731048960567,0.00453847549834263,0.00873545895223615,0.00318873197427805
"2554",0.00126891324123846,-0.00889773331518162,-0.00213046534719108,-0.0118130025310037,0.0111046730492896,0.00464072696773887,0.00500574219360517,-0.00212598014244547,0.00638973421238043,-0.00190709233946518
"2555",0.00156284588446454,0.00174563728176347,-0.00310560456499609,-0.00311862243565053,-0.00590114027821276,-0.00358247299555503,0.00522967960122633,-0.00399459922229684,-0.00484539694683539,-0.00254780134871879
"2556",-0.00269924537597099,-0.00174259534236676,-0.00253119263241841,-0.00964530310053924,0.00370998866038974,-0.000472721177697144,-0.00396390938048807,0,0.000923438526105436,0.00383143097049166
"2557",0.0139976126076811,0.0117208513778566,0.011711932645359,0.0155304035325612,-0.0167561098608832,-0.00696705592473612,-0.00310905399755845,0.000802054498062921,-0.00142585755030133,0.00445286527660071
"2558",-0.00629735372753171,-0.0036973925215037,-0.00945396507770557,-0.0176257193461409,-0.00359922799460299,-0.00286307980221256,-0.00411677093745944,-0.0125566710319954,-0.0124306738187582,-0.0158327854283856
"2559",0.000629381564045906,0.00841174127417554,0.000584232424516884,0.00765158312162728,0.00260410277387635,0.000957510829813435,-0.00237997397937695,0.00405833347214402,-0.000595339333299139,0.0051480673719293
"2560",-0.0029777352392526,-0.00515197933218881,-0.00233597423016452,0.000523773546083239,-0.00477570963343277,-0.000191436964855574,-0.00464613474526876,-0.00161686751653067,-0.00672284049488825,-0.00128045807361343
"2561",-0.00298703828645241,-0.00567208589159396,-0.00234144378250178,0.00104677419273358,-0.00303120773647392,-0.00143490764203147,-0.00428908098854786,-0.00485836235030701,-0.00805347834087144,-0.00448725015697193
"2562",-0.00185641960026983,-0.00421626074793802,-0.00312929310750232,-0.00941167710692248,-0.00540442604082569,-0.00335211393305734,-0.0153299637324174,-0.0086790846591186,-0.00621869931092334,-0.0225369177448197
"2563",0.00126820234268776,0.00797007402280592,0,-0.00791767631638118,-0.00798079254594364,-0.00278743400682369,-0.0127379481839037,0.000547385898523212,-0.0051277334456411,-0.00856391818071489
"2564",0.00350405748942473,0.00889542587552472,0.00725925545124384,0.011173212724702,0.00350894466170493,0.00212044202987438,-0.00247624363511667,0.000273365495677913,0.00218397831585593,-0.00930240351013967
"2565",0.000505003811898552,0.0039187624701662,0.00506413214011769,0.0139437810553684,-0.00631124404042438,-0.00250063349259066,0.00156784090784545,0.00191348776610245,0.000174311365286783,-0.00134129435353814
"2566",-0.00382671895928832,-0.00731890831984305,-0.00697660464156658,-0.00570837810110747,0.00480637128308392,0.00106075806648609,-0.000913334951957556,-0.00818538686360715,-0.00540347752141324,-0.00402956400638621
"2567",0.00865346807698697,0.0135169545735745,0.0101482766939005,0.0260959108673648,0.0122148966674109,0.00876399516743764,0.0184099194010034,0.0159559057780205,0.0186645368384717,0.00876603378785168
"2568",-0.0019669225702339,0.0104267189554459,-0.00193213992819286,0.00610375241894068,-0.00506338521723915,-0.00276837158540799,-0.00166683455732486,0.0119143193192062,0.00412905806451613,-0.00133694889041081
"2569",-0.00175610784859881,0.00191963418032004,0.00329092332896663,-0.00176939639504703,0.00627678805648557,0.0026805796077114,0.0042378373214973,0.00263636744525408,0.0022273193979101,0.00334674345417874
"2570",-0.00109690831120368,-0.00191595624522367,0.000192916551013722,0.0116485841285048,0.00429853146677805,0.00238703674289154,-0.000383724927288331,0.000804845497890838,0.00444485861090449,-0.000667102292611355
"2571",-0.0128396789882845,-0.00359978898565694,-0.00771610592965055,-0.0110138657863131,0.00830891702983849,0.00333405947462961,-0.0031980326324994,-0.00750668009223943,0.00876520281226778,-0.00534051833327187
"2572",0.0023532349836497,0,0.00136083816258492,0.00480895759237554,0.00399551315558,0.00189885030496661,0.00051336269804958,0.00270151796829343,0.00244643999960825,-0.000671062731966487
"2573",-0.00106701752946003,0.00120424723030488,0.000776582510718882,0.000251817771555141,-0.00140954953448558,-0.00104270531058959,0.00743970518262826,0.00404074167533519,-0.00134649497018424,-0.00201488568513231
"2574",-0.000726443133959309,0.00360844881822842,0.00620753347389047,0.00251840786784929,0.00356981049826244,0.000569317242158141,-0.000707065600293433,0.00295149963815078,0.00160110392855994,0.00336476113458128
"2575",-0.00102623015747316,0.00527311868793201,0.000578424903030283,-0.00276320337007108,0.00455023215144723,0.00246476037019483,-0.00681730068228059,-0.000535068511630099,0.00563686685481346,-0.00134129435353814
"2576",0.00727676540995481,0.00023843231029308,0.00847779050997111,0.00277085981926151,-0.00667047406185139,-0.00340448961907047,0.00440338644036253,-0.000802623440675609,-0.00409937257675375,0.00604431144893303
"2577",0.000934985710196568,-0.000953423816419052,-0.00133735785228317,0.00175828460679561,0.00596904385480701,0.00284689936425386,0.00438408163473891,0.00267848416424088,0.00243616429405091,0.00934580402420737
"2578",0.00318392838194725,-0.00381788187884613,-0.00554824950578392,-0.00526581051277752,-0.00807653698832289,-0.00283881753641424,0.00295296150330815,-0.00534334896973299,-0.0072069134801489,0.00396826774429404
"2579",-0.00232746763853919,0.00239530488338602,-0.009234243994378,-0.00705828412172327,0.00290806155675538,0.00199290727320367,0.00473631986764533,0.00456640668411112,0.00211023886122863,0.00197625751826047
"2580",-0.0017391526787599,-0.00382314715306309,0.00504856245789309,0.005585115599686,0.010086902427322,0.00492255179005419,0.00089190037153708,-0.00106972170578712,0.0053065784593449,-0.00394485458956617
"2581",0.000637283169812486,0.00143906781298697,-0.00347751898115156,0.0005051047989586,-0.00542476231351385,-0.00141587999260562,-0.000891105594126751,0.00214141985285354,0.0022622958066576,0.00990112731437764
"2582",-0.00297262366128581,-0.00670635680364251,-0.00697961417527004,-0.00302812469026936,0.00305747936702749,0.00189064053783583,0.00025479870902001,-0.00160263297956076,0,0.00196069013709699
"2583",0.00281121113330585,0.00337593631499433,-0.00507607934606946,-0.00177174407320924,-0.00148287509372325,-0.000660360747531952,0.00687823213873728,0.00909585024748027,-0.00367833965026731,0.00260929445926572
"2584",-0.00101941036347009,-0.00144214929942332,0.00215862008465884,-0.00177477996801234,-0.00404265224083677,-0.00302098874497392,0.00113857559032127,0,0.00234937909045141,0.00260250376062299
"2585",0.000595314018623005,-0.000962602424151027,-0.00234977849809492,-0.00406405470104532,0.00463897843333338,0.00179890058158505,0.00694951708394864,-0.00397671643991904,0,0.00778704458108392
"2586",-0.00118999131200481,0.00602260777388453,0.005102916886631,-0.00229531137595762,0.00948297571583567,0.0046316763272225,0.00552147786027746,0.0090497876290847,0.0144818601580603,0.00193185131067319
"2587",-0.00438170086903655,-0.00119730016460229,-0.00331953410031871,0.00485687223381781,0.00547277344458164,0.00310458970374206,-0.00224636373987896,0.00580334369110247,0.00684870852630226,0
"2588",-0.00649496884451228,-0.00695274391045941,-0.00842471471963524,-0.00432457389914864,0.00308741051721695,0.00300128913550224,-0.00200126180862059,-0.00209808298267922,0.00475332744025558,0.00321332361178372
"2589",0.00885999658218561,0.00627714605303065,0.0106696964283806,0.0104750972642398,-0.00307790775245098,-0.00158968491601219,0.0125329852510305,0.0113006938932059,-0.00293637851445971,-0.00576545622459146
"2590",-0.00298429909160014,-0.00527828451928669,-0.00312792601824285,-0.0126423033537344,0.0130800198695031,0.00571319604843312,0.00235188665138941,0.000519956198073768,0.00474478083679286,-0.00386605894290903
"2591",-0.0018385255204586,-0.00337682983485821,-0.000588407500659582,-0.00614568124507953,-0.00545292549275156,-0.00260750664927012,-0.00160557109828863,-0.00831180059958381,-0.00887475166910923,-0.0174644522676406
"2592",0.00813912711454079,0.00774458271198109,0.00608333701858621,0.0123678657302932,-0.00387053275130667,-0.00224089830845664,0.000618504758128191,0.00392895826744466,0.00188939451517145,-0.00394991328905014
"2593",-0.00318697453454775,0.000240254970751641,0.00370579830383289,0,0,0.000467993852801607,-0.0039555358899761,-0.00495737964158471,0.00286978519899783,-0.00991407848530956
"2594",0.0109979254532291,0.0362543990727437,0.0069956452875235,0.0142528805525413,-0.00493748561813045,-0.00205775673939024,-0.00868696321114237,0.00498207769210834,-0.00678599471483921,-0.00333780678179185
"2595",0.00581860997861749,0.00880449334264033,0.0036665275893617,0.00878303061256203,-0.0120395047130791,-0.0051551090812505,0.00287918956691136,0.00417420939639923,-0.0101251479224939,0.00468855149106728
"2596",-0.000628747296756105,-0.00390452220996029,0.00115365505637066,-0.00373135263953883,0.00551681979938312,0.00263789873436204,-0.00661582110796055,-0.00363731165268755,0.00490641164241157,-0.00533332912498308
"2597",0.000838793795045145,0.000691712010259637,0.000768331451396431,-0.0012484068936307,-0.000327631622622948,0.000657834439124816,0.00113099279588491,0.00130389816880783,-0.00372390776974207,-0.00536192604130525
"2598",-0.00217930642425623,-0.00115215708641392,-0.00479764387472803,0.00149989649507831,0.00221159344296984,0.00103289640771775,-0.00928833225982861,-0.00572941165631136,0.00315639175310567,-0.0026954503170562
"2599",0.0025201001899462,0.00392163608598328,0.0038565853640351,0.00574126001337727,-0.0083130043108971,-0.00216064850479114,0.00608138509797662,0,-0.00910821418667418,0.00202706893995463
"2600",0.000377233680258771,0.00689335437167027,0.00307333064143367,0.00719801280754484,0.00512048540917398,0.00207110509265851,-0.00251856396748429,0.0112625867988345,-0.000167092841432237,-0.0107889326307644
"2601",-0.00121478842466938,-0.00251025667206284,0.00248936617333029,-0.00665354066462209,0.000657440806270726,-0.00206682448194828,-0.0119936655813659,-0.0046619913918603,-0.0139573670880507,-0.00408999375384422
"2602",0.00117419071171576,0.0148707412700237,0.00248332510321436,-0.0111635113175481,-0.00492698525819635,-0.00226001820059629,-0.00434440680872195,-0.00208173503081199,-0.0100864720269586,-0.0239561487734999
"2603",0.00393715904546821,0.0114967950229403,0.00552590843140677,0.0082789976501676,0.000907709753131591,0.00018858049581727,0.0096253762701517,0.00573675962700704,0.00188373146773069,0.0140251252850372
"2604",-0.000166982580409147,-0.0104746457932766,0.000379139419816266,-0.000248747597336507,-0.00544147853111021,-0.00245255495952434,-0.0057200693290661,0,-0.00222204935950687,-0.00414932118355293
"2605",-0.000917856183288102,-0.000225221852377167,-0.00322039892211023,0.012692806670304,-0.0000829534957866862,-0.00113525451816554,-0.00536955069108824,-0.00103730263769186,-0.00599569164882219,-0.00486111622344032
"2606",0.00179569038708571,0.00270309889390408,-0.00456096508161852,0.00663544847801134,-0.00116067178434964,-0.000378436579475561,0.00539853841677496,0.00103837975174725,-0.0000861869861390474,0.0160502406843015
"2607",-0.00204266920328111,-0.00292040355568213,-0.00267273324085981,0.00219727141567994,0,0.000757692072218097,-0.00536955069108824,0.000518377045277019,0.00396414164112247,0.0041208935885988
"2608",-0.00167098827434642,0.00788621818787094,0.002488493427939,0.00414137165738016,0.0075529419319178,0.00511127947340206,-0.00269944557541957,0.00181386698891539,0.00283263519313293,0
"2609",0.00552334502452068,0.00581281152505864,0.00286425112387723,0.010189150448878,-0.00271829532202184,-0.000659408051852495,0.00360899835875661,0.00517325451344419,0.00265340233410249,0.00547195189069516
"2610",-0.000915411700343371,0.0102244380615419,0.00076158815866556,0.000960857668476978,0.00371711471554859,0.00131930658989976,-0.00565052659974108,0.000257314848325141,0.00435379037351713,0.00136059565705837
"2611",-0.0177441353430684,-0.0138613231578141,-0.00152215709143322,-0.0170346581617168,0.0145667435471653,0.00799925815552904,0.00529519914391496,-0.00360151140161591,0.0181895364523665,0.00679338516144568
"2612",0.00402859277772838,0.00133869235760731,0.00266772066206955,-0.0165977262744018,0.00113555846504165,-0.000280161985069971,0.00269783255771028,-0.00335656312506505,-0.00818100836312718,-0.00269901859172683
"2613",0.0065042304485039,0.0131461891803255,0.00817174907096829,0.0213453758787325,0.00234968866106078,-0.000279933498884333,0.00589351939440363,0.00595828666439657,0.00496594571106734,0.0196211203497609
"2614",0.00507724608151006,0.00241916512798546,-0.000565558928756871,0.000971986489439747,-0.00274827489905916,-0.00112124615600295,0.00292965545390067,0.00103014544421032,0.00418760461997314,0.00663567772410345
"2615",0.00221296460437159,-0.00153585800142664,0.00132036443976702,0.000971355048884126,-0.00672773857121467,-0.00261825879061683,0.00228600489424036,-0.00205792875612376,-0.00633864042804599,-0.00329593395865624
"2616",0.00233274509492465,0.00153822048967367,-0.00150690202328696,0.00388060941339075,0.00563069040318376,0.00206240135247082,0.00671579991958571,0.00386680839115816,0.00394495554763252,-0.00198416790706935
"2617",0.00477948629852976,-0.000877588658384054,0.00264104844718038,0.00483195880580767,0.000324604308653109,0.000561572525318077,0.00213961226679338,0.000256997499481493,-0.0010868489165885,-0.0218687617841493
"2618",-0.000206802582636501,-0.00483096524461157,0.000564356441123515,0.00360674870331823,0.00170367181638698,0.000654616762342242,-0.00615428071509805,0.00154029117873744,0.00887176074141882,0.00745254240077342
"2619",-0.000868820269268489,-0.00154457291633758,0.00206864685733166,-0.00527077086957162,0.0049399931467391,0.0025233962656499,-0.00391754133295907,0,-0.00331841709541714,-0.00806996786866232
"2620",-0.000248443363619066,0.00309390049654845,0,-0.00770701086025938,0.00249834356812206,0.000466256701494805,0.000253634407532344,0.00307617610336064,0.003995372099179,-0.0108473798076169
"2621",0.00795223313837257,0.00638914542359648,0.00900724155297561,0.00849502730933982,0.000104637793020945,-0.0005224996889448,0.00405877836077484,0.00920007659871658,0.000829033307186977,-0.00685405688185781
"2622",0.00332842252234089,0.00656737479486802,0.021015336472177,0.00505426763831496,0.0118405557562862,0.00438827061033065,0.00985368124998898,0.00734358953477776,0.00737243201315074,-0.0048309230214546
"2623",-0.000737171291897765,-0.00587207795883682,-0.00382510462257657,-0.00119749208412412,-0.00620934665421313,-0.00167351925889736,-0.00312753486301742,-0.00276526843412084,0.000986777395059812,-0.00554777457712019
"2624",-0.00319691091519936,-0.00371909064967268,0.000731350574751932,0.000479571116265065,0.00544718038517877,0.00316617623137905,-0.00501944393137388,-0.001512098611123,0.0112543741578648,0.00697340510093514
"2625",0.00185037388262499,-0.000219583880515017,-0.0003654080459915,-0.00119804473795015,-0.00478027994679242,-0.0018567020746123,0.00416207199959806,0.00403896286954275,-0.00528026816052429,-0.0138503695092584
"2626",0.000492347810953753,-0.00373376981907603,-0.00237606852510197,0.00599782048993647,-0.00264159353578786,-0.00158076615887048,-0.00163288596318623,-0.00402271527192455,-0.0065332382164125,0
"2627",-0.00151780126918188,-0.00286613471300101,-0.00897776394559013,-0.00763154870963623,-0.00152491610496286,-0.000931432131144216,0.00641614682365366,-0.00732166623391062,-0.00912454567818255,0.00561797306157019
"2628",-0.000205335812921148,-0.00508499660352491,0.00314298083347109,-0.00528723774775308,-0.000321594088146804,-0.00018632387496087,0.0066248200170167,0.000254513785849397,-0.00149328022653661,-0.0090782320655145
"2629",0.00488994912190788,0.00577764262029734,0.00552892691490992,0.00483195880580767,0.000160917613847511,0.0003728751688854,0.00211113604532964,0.00991589105887836,0.000997025581613187,0.00422841721504996
"2630",-0.00126774623981007,-0.00176753891338044,-0.000549829488926901,-0.000240477415349605,0.0154364509784344,0.00521988572713528,0.00322176699747523,0.00251758357903986,-0.00547811241339369,-0.0175439077995795
"2631",-0.00192428340029038,-0.00996020442049483,-0.00971943481584525,-0.0103414687737421,-0.00158352677993834,-0.00176161235581662,0.00345835068727585,-0.0050226406106324,-0.00417292605575026,0.00428580271427803
"2632",0.000218486666245576,0.0111782095723296,0.00407403975198628,0.00170113270823391,0.00198234846031475,0.000557251361201772,-0.000615319383985957,0.00349120789907342,0.000167582970164393,0.00426729339038379
"2633",0.00832523503787064,0.00375872868494964,0.00313538684817538,0.00994651446528771,-0.00142444948430542,-0.00278553076391286,0.00172427683985088,-0.00126962591253721,-0.00762523906905432,-0.00637392368741607
"2634",-0.00674416515847009,-0.0104541852176463,0.00033313477758834,-0.011052620909646,0.00895616634475638,0.00251398440049755,-0.00331987622632457,-0.0162726109089109,-0.00211095161698893,-0.00997862781066583
"2635",-0.000247017724704257,0.000226743735882273,-0.00147987635983204,0.00219630612481714,0.00204255667427722,-0.0000927248131284975,-0.00394772860063608,-0.00258471753559442,0.00287694195295307,-0.010799137029343
"2636",-0.000452655397962687,-0.000906550664983463,0.00203786751070578,0.00511314565961385,0.00219481251118725,0.000928681358615568,0.00198178943157923,-0.00414609603310312,0.00337496633584977,0.00145565913800816
"2637",0.00119429845411911,0.00340300837603924,-0.000739595308469787,0.00532946385358346,-0.000469285175990208,0.000278315456205824,0.00395553588997632,0.00442374176639571,0.00428861426654237,0.00436033063266361
"2638",0.000658012028253996,0.00339127329111566,-0.00277515856083066,0.00963860330116684,0.00375654655797719,0.000834861385007546,0.00640229411045135,-0.00207275189649625,-0.00895921460269622,0.00217088652750053
"2639",-0.00805619390485157,0.00247854770355893,-0.00241185774635211,-0.0116945671781526,-0.0106814688786249,-0.00491245531889961,-0.00591208787017683,-0.00519197787236914,0.00380193474314017,0.0115524115461247
"2640",0.00895038837195083,0.0074175000309622,0.00446335989229851,0.00772764660200442,-0.00331009602691579,-0.000931432131144216,0.00136563855882432,0.00104388795535781,0.000757545673891968,0.00642396808240298
"2641",-0.00878876814201657,-0.0111557491812805,-0.00999805134243037,-0.0127005622180066,-0.00838134433443116,-0.00372929086633644,-0.0109113962511117,-0.00469255172819449,-0.00487806551929248,0.00425518775965816
"2642",0.00186440600263404,0,0.00336637967379771,0.00461167059476519,-0.00231232784909408,-0.00233928759051483,0,-0.00209530972812044,-0.00253552231237308,0.0204803110442378
"2643",0.00169554379090631,0.000451169342021274,-0.00484619307602763,0.00579843764276089,-0.00321968982279963,-0.00367299155387835,0.0106558898304976,-0.00892411580296615,-0.0163531693701027,0.0103806233302839
"2644",0.00231215390095008,0,0.000187215505753402,-0.00192169550406418,0.000241114224354355,0.00075396937658434,-0.0112876531034896,-0.00158876162276589,0.00370403148260934,-0.015068498558463
"2645",-0.00914462535319804,-0.00360852486771113,-0.00730345909690511,-0.0120337541608667,-0.0082737145546089,-0.00188427529583812,-0.0174381026422691,-0.0050399747908616,-0.000429076564428699,0.000695472358283933
"2646",0.00648525054821847,0.00203714481477402,-0.000565810604726713,0.00194884747945867,-0.00599358662512595,-0.00160446301684058,0.00485160582921207,-0.00106605777811564,-0.0102172404033893,-0.00972898790088284
"2647",0.00107376684064842,0.00225897595398572,-0.0026424040852695,0.0094821749011238,0.00146674427899862,0.0013235764351498,-0.00736973842788524,0.00186808144093131,0.00164817836266629,0.00421046853524154
"2648",-0.000742611973443719,0.00135222438483185,0.0068129134632644,0.00818877291389941,0.00170837103195987,0.00132189677288208,-0.0011519538556618,-0.00612678511174625,0.00129905602061964,0.00978337842656662
"2649",0.00751487727509548,0.00855287671231553,0.00695479401550037,0.019350187457204,0.00690449084197731,0.00292295015930222,0.0125592326097224,0.0069684064851776,0.00354606460267948,-0.00484429563586741
"2650",0.00168018719893914,0.00423996933645299,-0.00130661196789217,0.00492161797262192,-0.00629260118215691,-0.00103411332446279,0.000379907105910071,0.00452500494185948,-0.00180986815314899,-0.000695400785539535
"2651",0.00466401367348612,0.00622230573685134,0.00242987082172164,0.012593256101108,0.00121812472982374,0.00141164867675658,0.0101212273216698,0.0135135868834237,0.00820235710585404,0.0111342268915033
"2652",-0.000121995673945663,-0.00154595701699711,-0.00130520848532278,-0.0046061951207832,0.00275673228072626,0.00122195993299323,0.00400825286247319,-0.00235305404548869,0.00445323296531375,-0.00344110942841314
"2653",0.000529373076654016,-0.000884883610975717,0.00522777406657493,0.00300786443131829,0.00873283007383829,0.00366081025087994,-0.00249515681958135,0.00943401925300336,0.00699121828807892,0.00414366093869045
"2654",0.00541404139157486,0.00199252008747086,0.00408619732501592,0.00830455444909739,0.000400757324678258,0,0.00800397077744242,0.00700941040889069,-0.000253992039166984,0.00894087224434292
"2655",0.000445319215181872,0.00552363757864138,0.00369956538323235,-0.00114401852348367,0.00288474352046419,0.000280485429446475,-0.00397036319965838,0.0043826562999445,0.00135497965184661,-0.00136337802319941
"2656",-0.000890237744159306,-0.00593259612023034,0.00184298376289238,-0.000687040818165063,0.00423451772056893,0.00177687506859781,0.00211774762446271,-0.000256692441097828,0.00862655630288489,-0.0136518315761254
"2657",-0.000243013854036911,-0.00309483718231918,-0.00202354508283809,0.00297952545029267,-0.00389857470945143,-0.000653325903290591,-0.00261030195673995,0.000256758349025166,0.000419218507140329,0.00207609617564697
"2658",0.00243086521421731,0.00221737917276554,-0.00350228380531203,-0.00251362868035343,-0.0130189824644729,-0.00560390197970406,0.00124629406435384,-0.0015401546465873,-0.00326879562934856,0.0110497861959944
"2659",0.0000404259233230952,0.00774339559958115,0.00332956250041172,0.00824738037952089,0.00161852695949549,0.00319323959742213,0.00535212838185051,0.00437017353197433,0.00807264561171617,0.00956278073642225
"2660",-0.000929606057609167,-0.00461030944993279,0.00331862877971778,-0.00545334299985967,-0.00492852250178288,-0.00159153268857137,0.00086658165147413,0.00179157976284583,-0.000750717402837386,0.0060892964033703
"2661",-0.00117316607847007,0.00110279713452899,0.00294003911957152,-0.00045694114894046,0.00592727524631975,0.00168793589957916,-0.0021027543991099,0.00383265017338208,0.00751315629423854,0.005379955507687
"2662",-0.00056692384595558,0.00264367474048122,0.00329797491808526,0.0011428750990119,0.00121054860089642,0.000280896432650835,-0.000123894953048875,0.00152680382852455,0.000497124857119502,0.00602005367344782
"2663",0.00222870431881095,0.00483422456970706,0.00584372181839021,0.00296805874005535,0.0070212058831951,0.00248383179166178,0.00446313155845468,0.00330384057894473,-0.000828140786749532,-0.011303174426881
"2664",0.000485358150433601,0.00109327485468547,-0.000544773836603452,0.000910432279300988,0.000561623398552591,-0.000935255952501435,-0.00629478429376784,-0.00253287918521317,-0.0020721093730276,0.00201745736003356
"2665",-0.00193997790923439,0.00152907250372425,0.00254317691005546,-0.00409361919403362,0.0103440231960659,0.00346286746484781,-0.00347762868839052,0.00126965547653568,0.00157802322960099,-0.0073824498756202
"2666",0.00182211766448548,0.00196296891110181,-0.000905963959782596,0.00365390834205082,-0.00849209747505575,-0.00270467144862796,0.00336519039493677,-0.00202909128917772,-0.00779495838112476,0.00202830017005384
"2667",0.00185916332618596,0.00108837067232814,-0.00036268011231666,0.00682577784843352,0.00112069058682773,0.000561335598459056,0.000745236883027411,-0.00355769312416709,-0.00117007937868652,0.00202433339157682
"2668",-0.00246085746668567,-0.00652314776581264,-0.0010884729684264,0.000225992260157071,-0.00359810938970628,-0.000841185693946978,-0.00546159048893513,-0.00382559977756991,0.00292861680313594,0.000673322171594659
"2669",-0.0000403842195622062,-0.0013132520322876,-0.00617514530841046,-0.00903735857784704,0.00545657402574218,0.00121602505478102,-0.0017474275021353,0,0.0120974218913947,0.00672959153000807
"2670",-0.0141153786124706,-0.0149024915623966,-0.0104166062552177,-0.0237119124979532,0.00853954029927251,0.00373717208366631,-0.00762698208804502,-0.00972853699814558,0.00741901751576979,-0.015374396255745
"2671",0.00147701279973944,-0.00200217660450175,-0.00147741668438484,0.0023352693497698,0.000474736225117178,0.00111707260044325,-0.00478751959032653,0,0.00474594554247565,0.00339445675241579
"2672",0.00991302166277697,0.00735612993224066,0.00739782030394753,0.0102517679627521,-0.0051413023725202,-0.00241757750361948,0.0153181869797578,0.00672171437307023,-0.00708529190418361,-0.00879568904694039
"2673",-0.00012157879742003,-0.00110645775601792,-0.00128509955099232,0.00115315458489529,-0.00421356438080611,-0.00298228825815849,-0.00286776229249186,-0.00487924368194959,-0.00770993286925747,-0.00477816212774163
"2674",0.00174429777905405,0.00531694187724674,0.00330873352210448,0.0103663142193597,0.00367270962999333,0.00186963878652846,0.00437666118839686,0.00851618735377824,0.00735658768333813,-0.00274344684758798
"2675",-0.0155907687137479,-0.0125605406702601,-0.0067790070293885,-0.0127680483545705,0.00747756574725966,0.0035456264313336,-0.00684778964342736,-0.00639721905064461,0.0050873470479853,0.00275099405355195
"2676",-0.00156324177917044,0.00066936559595776,0.00442728699882,0.00854507063859167,-0.000236994772004895,0.000186160779940936,-0.00739616276940258,0.00386312812186063,-0.0015511062380783,0.0178326868731391
"2677",0.000782712871222335,0.000892113592482202,-0.00220384791861916,0.00366387559399284,0.00244839035443722,0.000650523926853941,0.00896689727191324,-0.000256590609398866,0.0037612345765845,-0.0121294223954782
"2678",0.0104571973357963,0.0057930921149274,0.00202460472124288,0.0111795865948021,-0.00386051184131297,-0.00195099934288712,-0.000876018172116688,0.00179620687974946,-0.00448031110328595,0.00272854600406491
"2679",-0.00358549597364732,-0.000221498675187615,0.000367420217837644,0.00473819682208965,0.00680181402945745,0.00344431864830508,0.00826842300717234,-0.000768469564635943,0.00376400461307602,0.00884355670473025
"2680",-0.00233070178157235,-0.00132945275996066,-0.00514139955757087,0.00314397336631611,-0.00369205099507997,-0.00157694880221326,-0.000994094458116712,-0.00358890950739599,-0.00309771750383503,-0.00067436901525264
"2681",0.00233614664271453,0.00710010734645317,0.00332224588584795,0.00582040916624837,0.00386316894271399,0.00167207308797157,0.00472640382214307,-0.00128619462866519,0.00367975301594758,-0.00202419449601332
"2682",0.0000409630100031144,0.000220373144092623,0.0011037483717955,-0.00356093731937857,-0.000628208507072125,0.000927717192391819,-0.0050754430429395,0.00309108845577177,0.0158872741712119,0.000676053664256049
"2683",0.00114476031083277,-0.00396475647143568,-0.00202139079060126,-0.00178701026281025,0.00322231057836997,0.00231674714661145,-0.00149318249651342,-0.00205441524523564,-0.0021654021627171,0
"2684",0.0047375832453842,-0.00176930462831459,-0.000552420750399518,0.00156625109829589,-0.000313417395879312,-0.000832164447078232,0.00535845669570589,-0.00154390851797515,-0.000482213478254612,-0.00743240066882345
"2685",0.00601606246075392,0.00731078617567094,0.0079219264592747,0.00156399256353579,0.00297787265380478,0.00157323392492237,0.00644488032303414,0.0108247011258826,0.0117401012243479,0.0279101820157066
"2686",0.00141421050328305,0.00219905243840413,-0.00402106618215214,0.00736118616300607,-0.00764906975543722,-0.00294264452435766,0.000123287293481766,-0.00382459460027484,0.00190747099030353,0.00132448516535044
"2687",-0.00718207122247283,-0.0063636964782201,-0.00440453674104513,-0.0130648161361986,0.0158578671252576,0.0069601622833475,-0.00209318724658858,-0.00102361087160507,0.0111058307330769,0.00198403176737982
"2688",0.00341360874162211,0.00706698856664167,0.00423964013301248,0.00650674559192788,-0.00613542787873189,-0.00239585649416985,0.00197404720141603,0.00614891287812136,-0.00509964698807197,0.00990112731437764
"2689",-0.000121269858061379,0.0089912922443971,0.00587365977921239,0.00735616813996631,0.0102367606889668,0.00434153519233127,0.00652740629234438,0.00814884170789609,0.01040932908145,-0.000653653071059468
"2690",-0.00117473845851435,0.000217403556616036,0.00310226013536963,-0.00663867043776079,-0.00216578204374185,-0.000735808200046595,-0.000611826458065678,0.000505391776847164,-0.00124876292637321,-0.0111183607233376
"2691",0.0106658082957851,0.00760530424850847,0.00454791071242133,0.0133660738347574,-0.0119380636621491,-0.00570702548464541,0.00844751887817385,-0.000252950342726321,-0.0139095021183909,0.00198403176737982
"2692",0.00337071792930632,0.00452875859730373,0.000724252617180454,-0.00109915992224308,-0.0052563670457717,-0.00240710537375055,-0.0100764646969405,-0.00429271789676933,0.00293205479147218,0.00264029608816352
"2693",0.000479933252762521,-0.00601115256179829,-0.00199043743718785,-0.00528153824431399,-0.00394354122700147,-0.00204120849261369,-0.00367903268012681,-0.00735493551853128,-0.00750629752696419,0.00460829992672163
"2694",-0.000319906824606142,0.00323984068423622,0.000181297698183647,0.00265471965681052,0.00411751981423358,0.000185820998266806,0.00615451055709748,0.002044036466053,0.00437865612309007,0.000655366512221311
"2695",0.00134633336678558,0.000430596043653697,0.00145038363402228,0.00595765753177235,0.000394177038070431,0.00120870472009549,0.00415942935586888,0.00324043119624329,-0.0049936983197939,0.00458415661069123
"2696",0.00212688831287156,0.00193668671828173,0.000180926721635277,0.0035096434422246,-0.00575442389013625,-0.00390047622407552,-0.00536064872327879,-0.00281989453748865,-0.00932046530168462,-0.00130376311982083
"2697",0.00100108792064235,0.00472511299926537,0.00579189538606006,0.00218561644096082,-0.00245774148561717,-0.00111847956896072,-0.00771662835142217,-0.00308492083893019,0.00209072047209125,-0.00195826488688433
"2698",0.000359988310639769,-0.00299277192873426,0.000359873684092626,-0.00458008517888031,0.000715387199296424,-0.00195954569632262,-0.00246898985488819,-0.00257850424966122,-0.00802439396506838,0.00850230752397341
"2699",-0.00267930703672647,0.000857660845482888,-0.00395756201245245,0,-0.000555973209028893,-0.00130932623626989,-0.00321725007868023,-0.00698026669289498,-0.00760397166468274,-0.00389106408858941
"2700",0.000200492568461552,0.0021422573226173,0.00108376585898862,-0.00569677646657951,0.00286062904971596,0.001778927683173,-0.00595908539540779,0.00442596111890414,0.0045647049233779,0.0039062636106455
"2701",-0.00204463769740693,-0.00769566323515347,0.00216480850546685,-0.0169678115838858,0.00625994587851153,0.00299106080556721,0.00537028459464528,-0.00544331426267519,0.0104673890046638,0.0168611887231829
"2702",0.000602660484037232,-0.00301591263000622,0,-0.00268990241360501,-0.00181127765409073,-0.000838856084123818,0.000275425971241861,-0.00208488106557636,-0.0111619690930858,-0.00892858080554015
"2703",0.00389425497181928,0.00172859523696456,0.00198014000568913,-0.00359634595531921,-0.0150677447754115,-0.00512965045745539,-0.00801601554629727,-0.00444004285669763,-0.00942013975491429,-0.00386108364400783
"2704",0.00119985542637346,0.00345122470334536,0.000718733637917746,-0.000676825436848105,-0.00296337901713783,-0.000187336606640165,0.0074496748557793,-0.000262099791770387,0.00188552217038396,0
"2705",0.00351492863496539,0.00752374686926305,0.000179451278659259,0.01151247600925,0.00224916697843636,-0.00121893899344594,0.00112788779228179,0.00708478888696273,-0.005155036454914,-0.00516788856168493
"2706",0.00433878296775325,-0.00192022717126594,0,0.00022314415014435,-0.00183116563982511,-0.0011376049937265,-0.00200284482295954,-0.00234499261387322,-0.00666232099584918,-0.00844151018349193
"2707",0.0021401399069918,0.00320648242649346,0.00592362169980376,0.0158410575511312,0.000965600127203814,0.00141189915221163,0.000752540266587998,0.00470085833372691,0.000496853535568054,0.000654869887072751
"2708",0.00118639768679452,-0.00170465343639781,0.0001783625295253,-0.000219568541018345,0.0000803215146958358,-0.000282120193747848,0.00639252591830264,-0.00519883407809918,0.00281383757653186,0.00130894998339981
"2709",0.00592515282358685,-0.0012806445795881,-0.000535197036823143,0.00746929128784579,-0.00377766572435445,-0.00103404326720036,0.00311379035204529,-0.00130656866235479,-0.0053643724579413,0.0111110931727056
"2710",-0.00113886779089012,-0.00085500292294205,-0.000535483626073141,-0.00501529585520832,-0.00282414416688603,-0.00122359344675405,-0.00360077293232897,-0.00183152882373239,0.00472949729661876,-0.0155139513659167
"2711",-0.00165112578046367,-0.00042774117279365,0.00125021201212938,-0.000657449123599219,0.00315558584412368,0.0011308164358399,0.00199381214489258,0.000262135712596034,0.00817578687507758,0.000656522276818006
"2712",0.00263833120198886,0.0106997799656545,0.00713514021220618,0.00986845878127807,0.00161331913767038,0.000376460211067187,0.00136782290267523,0.00707559768309052,0.00262123193608743,0.0118111334310549
"2713",0.001571015476999,0.00254070440467302,0.0051364396301985,0.00456028557673838,0.00193255867865005,0.00112925270427833,0.00422274646276621,0.00572487667284172,0.00318626628780616,0.00194549867153038
"2714",-0.00149018528364164,-0.00190069352877853,-0.00123346911334854,-0.000432437999934199,0.00425985351232061,0.000939774722519937,0.00655449927123763,0.000517100728653741,0.00081438227205477,-0.00129448070386373
"2715",0.00121756326152367,0.00169284116070778,0.0123499612189721,0.00908309543224117,0.00720295978778784,0.00338040388351546,0.00221152341989095,0.00284453920736349,0.00756775170939661,0.00972125587305173
"2716",0.00133344688808101,-0.00253498176100242,0.00453122015507978,-0.000642867565873062,-0.000715180237723545,-0.00168450762563832,-0.00502627777959042,-0.00128914795005619,-0.00686479567113552,0.0025674912770961
"2717",0.000705165181145162,-0.00381201147642141,-0.0010409396666472,-0.00514700425751702,0.00127229272873031,-0.000375282357058859,0.00086251474089627,-0.00103272112449659,-0.00683096684694662,-0.00128045807361343
"2718",0.000978617200084742,0.00425188500683493,-0.00104187931328936,0.00237119188118551,-0.00659170579191837,-0.00253152119308631,-0.00110798617287655,0.00439369164521053,-0.00376647024727261,-0.000641082861988718
"2719",0.000273681097441525,-0.00169364851738529,-0.00226021329151105,-0.00881722796603135,0.00175888742789598,0.00103394577553018,-0.000739383709166153,-0.0012866127785931,0.00591765440811454,-0.00448993064839287
"2720",0.00516044857352038,-0.0029685665544138,0.00226533342823521,0.00368853998474616,-0.0106137964413938,-0.00413211426732452,-0.00320699216578924,-0.00438022603260668,-0.00637305340610395,0.0051545684159735
"2721",-0.00388943935287756,-0.00319004766593245,0.00243382316750651,-0.00799839558164739,0.00177462622706037,0.000942816371767963,-0.00470161247263601,-0.00879920275064283,0.00156238794866881,0
"2722",0.00175711172158,-0.000640129090717756,0.00832464660729215,0,-0.00619951799727458,-0.00301482699704902,-0.00497276331533314,0.0015666241872212,-0.00385879300840419,0.0102564681117521
"2723",-0.00495013250466847,-0.00106738973649345,-0.00808399886624289,-0.0021789722318154,-0.00478017436812084,-0.00160643059974341,-0.00387295370481511,-0.00782074821382917,0.000164806722742883,0.00126895282363715
"2724",0.00129268496459289,-0.00235097738250478,0.00537538470984633,-0.00677014270075915,-0.00333785453532387,-0.00132500878243813,-0.00614579618010214,-0.00157650314903346,-0.00840540598937634,0.00443606490635928
"2725",0.0081761916249794,-0.0017138747520421,0.00758885418931698,0.0145117491637965,0.00661618355404348,0.00322201104768172,0.00454316540136568,0.00447383721345251,0.00473697324462785,0.00504724945748625
"2726",-0.00372498019924472,0.00579410551849846,-0.000342263778087104,-0.00628515641825811,0.00957470201635924,0.00359019647795766,0.00213552505218084,0.00104799332230843,0.00190235728862942,0.00251101593966951
"2727",0.00155767322246869,0.00512050667996933,0.00428079879334042,0.00937836942142067,0.000321490331252949,-0.000658812976897738,0.00188056419847138,0.00680440226852896,-0.00379756469406989,0.00250479097826695
"2728",0.0013222217707114,-0.000849104243377696,0.0056265404344451,0.00518593040109949,0.00445247634360535,0.000603809376310993,0.000750765131016129,-0.00441902846902553,0.00364633303466189,0.000624536740310377
"2729",0.000388500879768605,0.00254940917917112,0.00118683243441087,0.00128978808323366,0.00440891016032707,0.00132003719906693,0.00625150270022368,0.00391648512495091,0.000660564770369465,0.0062422403245177
"2730",0.00333867322693604,-0.00254292621972463,0.00237090410109864,-0.00515236920303475,0.00271362469730563,0.00160063372295594,-0.000621279825986032,0.0013003319905236,-0.00470335003377598,0.00620332494232834
"2731",0.00154767375310572,0.00212448487493355,-0.000168799818300647,0.011221374931971,0.00374069294229673,0.00122228110396749,0.0115628169284008,0.000259842591213699,0.00853920555780463,0.0191123283471131
"2732",-0.000695402371721943,-0.00826791229300139,0.00794179266743211,-0.00640198939252756,0.00420266211709275,0.000375335918987307,0.00712888550454527,-0.0025967318273431,-0.00361695842799903,-0.00604964843524292
"2733",0.00170080927922633,0.000641177324395059,0.00620281919344245,0.00472493032316446,-0.0022109849967471,-0.0012198772167149,0.00671229565956954,0.00937258465647584,0.00346504416685955,-0.00182590324516907
"2734",-0.00362766083421451,-0.00704957631778391,-0.00833051165773502,-0.00619909987092115,-0.00284879532595916,-0.000376107605841614,-0.000363792016166542,-0.00232149295314232,0.00411082802213669,0.00182924326638534
"2735",-0.000309946481561019,-0.00150604410324462,-0.00739248422147565,-0.00430209055276021,-0.0150796919508792,-0.00507664635883653,0.000606374966061418,-0.00180965787878118,-0.00818799659841141,-0.00182590324516907
"2736",0.000930058994298211,-0.00452487778485189,-0.00440085365245357,-0.00216030466408501,0.00209516314749392,-0.000472636712428032,0.00363600576507972,-0.00492108979847627,0.00148601506198331,-0.00304873877730882
"2737",-0.00232261733057137,0.00216432874287342,-0.00527028932008733,-0.00671135309887894,0.00675475884806653,0.00141827265538552,-0.00156999727060647,0.000780910606720697,0.0020608359090073,-0.0134557875869372
"2738",-0.00500519828790735,-0.00453560562476585,-0.00734918920091643,-0.00523107286220958,0.010862685268094,0.00358716979028295,-0.00858713324973659,-0.00130021191184682,-0.00123390920095268,-0.00123984494504614
"2739",0.00850095217885416,0.00650911151876765,0.0154958059377404,0.0208150971089545,-0.0086915174099419,-0.00253967689766621,0.0067096277131915,0.00937478367091971,-0.0000823820086522931,-0.00310368377575998
"2740",-0.00293882324083883,-0.00129334331546327,-0.00491690757008123,0.00493659868213348,0.00741257715555532,0.00132043494847944,-0.00460475375530678,-0.000258099575334403,0.0120263507079679,0.0161893255167598
"2741",0.00170640311853809,0,0.00494120300855938,0.00512604967877905,-0.000395580223472414,-0.00160116276467881,-0.00206968529317764,0.00258061952502664,-0.0126160099901025,-0.0079657033931777
"2742",0.00654278706996436,0.00539588224975884,0.00915575160183879,0.0133871489294548,0.00316619592209055,0.000188684100529191,0.00719762480618757,0.00592039979997638,0.0016487017005804,0.0067942881877463
"2743",-0.000884430768348432,0.00364966779358311,0.000671999375899235,0.00251633513994087,0.00323480785376051,0.00320655879566401,-0.00278591486353508,0.00230284163238048,0.00921730706580015,0.00552146022906941
"2744",0.00230964609515749,0.00919794861258705,0.00822695931452633,-0.00209171234248029,-0.00275242707246826,-0.00084625920347503,0.00206500112290131,0.00459536668459504,-0.00252790514216528,0.00305072465542766
"2745",-0.000499260162471815,-0.00635864007889553,-0.00432962699266826,-0.0146719615148461,-0.00141970928962754,0.000658761280818432,-0.00412120367936575,-0.00101644960535729,0.00416940810987576,-0.0018248551037251
"2746",0.0101447996196418,0.00639933112224766,0.00301040246727946,0.00744536427329523,0.00134247939168919,0.000188090776940708,-0.00219079705045777,0.00432448243966843,-0.000162859233691082,-0.004265696046719
"2747",-0.000608622973302997,-0.00402716446741369,-0.00200092303428356,-0.01583623786513,-0.00985877417462,-0.00319630964087136,-0.00121994260394098,-0.00658563521438738,-0.00626982340639715,-0.00673198010526599
"2748",0.00875497698502259,0.00106395962802708,0.0010024324930038,-0.010941892209768,-0.00334540597065125,-0.0031123386043157,0.00109929600127545,0.00484446320658916,-0.00770241717713527,-0.00431300522668032
"2749",-0.00207539278372681,-0.00361379574507503,-0.00450677732053417,-0.00563986297791874,0.0134944833361308,0.00369524572429181,0.0018299858084827,0,0.00404622632611429,0.00866337563776698
"2750",-0.00120999055229842,-0.00149360404960097,-0.0105633215462881,0.00196345140593968,0.000474056863773553,-0.000472000704836439,-0.00767199025720278,-0.00380617605993028,-0.00337195504143284,-0.0122698975885782
"2751",-0.00359668133342306,-0.00363239660731685,0.00254189659012449,-0.000653270989964483,0.00497591050179369,0.000755589462345441,-0.00589012894545426,0.00382071838678577,-0.00709688067337855,0
"2752",0.000190043470778667,-0.00171571248115487,-0.00371867313053231,-0.0135075811856634,0.00345798884482496,0.00207634179798633,-0.000370238517528931,0.00177622525743937,-0.00207779255319152,-0.0167702126206949
"2753",0.00315310809254665,0.00257788818493476,0.00644719705161889,0.00287085745191384,-0.00783199167789994,-0.00178963242272001,0.00407507794880635,0.000759856247711133,-0.0131590072457732,0.00315851657128929
"2754",0.00545295910410504,0.00514254249910495,0.0047201021933565,0.0116714813340002,0.0000789909706095937,-0.000754726178185283,0.00332060841427251,0.00379654259437134,-0.000084353111390878,0.0050378444325565
"2755",0.00301315533807633,0.0019185898783729,0.00335580261891066,0.00500665559058922,-0.0020523433350822,-0.000660904006159813,0.00110303424472269,-0.0017649121940031,-0.00396692258692799,0.00250629588749507
"2756",0.00176473412488165,0.000425465916426004,0.00183941102118457,-0.00671435223189976,-0.000395418184782614,-0.000850488288749895,0.00404064989456088,0.00303115462862458,0.00118634012056029,-0.00875007309041997
"2757",-0.000112398559400484,0.00212676683973667,0.00400613270487082,0.011993070450075,0.00751728893161308,0.00406646523731347,0.00207332464638377,0.00956936825502419,0.0086330595237738,-0.00441362391405054
"2758",-0.0040862816888616,-0.00594226374459028,-0.00465517803624971,-0.00732612172945091,0.00424079805803701,-0.000376875498849238,-0.000608409921110997,0.000249306676089578,-0.00201391293134034,0.003166583158283
"2759",0.00832753981404522,-0.00106738973649345,0.000501118606927919,0.00217071359304644,0.00375391661487767,-0.000188325914686871,0.00414007656436088,-0.000727008810516683,0.00210207685192976,0
"2760",0.00634126457286932,0.0132506551761458,0.0120200558964074,0.011262600189287,-0.00911592755412649,-0.00226164176897126,0.0055784953106579,0.00978438445401908,0.00461489343849641,0.00441919659547785
"2761",-0.00384049283305721,-0.00105464715164316,-0.0101459359118562,-0.00528343029170353,-0.0129735604865129,-0.00453339803925279,-0.0192564649320616,-0.0032300875097776,0.000751666230226267,0.00754251726589228
"2762",-0.000523851371167838,-0.00401185861603803,0.00134195712626428,0.00131145256333309,-0.0110732323615021,-0.00294127285607659,-0.0104388153749211,-0.00174465434525894,0.00267066432982821,0.0056144599261303
"2763",0.00205948333219386,0.00420375934602113,0.000670192274732306,0.0065488581569304,0.00582832179781323,0.000705058928102131,-0.00364176995113752,0.000749114071553203,0.00141500750303813,0.000620211184653829
"2764",-0.000261466158084755,0.000849928314172743,0.00468770042386457,0.00845802421419029,0.00136432854811663,0.000381055013856102,0.0063018325617199,-0.000498863662829918,0.00523650578067514,0.00433987205688369
"2765",-0.00119632946520987,0,0.000499959562221264,-0.000860230186418787,0.00296548857829593,0.000380899892951536,0.00488504747807461,0.00149745260228329,0.00686286577041728,0.0148148021084444
"2766",0.000486693460609811,0.00148620190855753,-0.00133248442615108,0.00258291245852194,0.0130254142524815,0.0042827843800024,0.00361432139527129,0.00648065167112555,0.00377766289999992,0.00243299406141095
"2767",0.00205725307689475,0.00233194272031767,-0.00233479041107731,0.00686984130997037,-0.000867532782373948,-0.00123201732980271,0.00583715979625476,0.0034672109474434,0.00507236345236772,0.00485430284159838
"2768",-0.0037703501191948,-0.000422941732748372,0.00183884562288483,0.00469086937655017,0.00157890704553965,0.0016128376910598,0.000247068609048107,-0.000740339836018511,0.0065120391780551,0.00301940706457482
"2769",0.00715733504954552,0.0067711028400963,0.00600693450716516,0.0188879207616086,-0.0107994207937171,-0.00331548616059352,-0.00506110561700246,0.00592719183296997,0.0121310147653697,0.00481637198410567
"2770",0.00632495906756336,0.00273221254936207,0.0137668161689519,0.00958144022710417,0.0047813302984463,0.00104551346279158,-0.00161288869981946,0.00564706971485895,-0.00263685173572759,0.00599165342118746
"2771",0.00421477843014473,0.0121567735683563,0.0122708915232557,0.0049514512350699,-0.000158578559307343,-0.000474634877408509,-0.0156581699996684,-0.00146485808071339,0.0051273754206056,-0.00119116894609306
"2772",0.00666398884758101,0.0068337265985785,0.00274782632482529,0.00862248144273225,-0.00285556949992161,-0.00123486355548774,0.00100999771596921,0.00440096496762399,-0.00103616292871167,-0.00357789130999808
"2773",0.00182882956802577,-0.00267376955682597,0.00580270346855039,0,-0.000636365878667777,-0.000475666558101384,0.00567543758982914,0.000243304072093942,-0.000159610625395157,-0.000598312713800175
"2774",0.00226320893723808,0.00144362073293092,0.000640936515176715,-0.00162836156945989,-0.013372478486519,-0.00475726465590287,-0.0115374512740504,0.00146022380206423,-0.00462848144008432,0.00658673582176394
"2775",-0.00152948350342907,-0.00329500427364937,0.00640618986660857,-0.00632012833265827,-0.00121009844205577,-0.000286766412597395,-0.0121797642544577,-0.00680421851614743,0.00240516309456029,0.00356925525226215
"2776",0.00729582518206273,0.00702486105650957,0.00668357020198562,0.00615517407671806,0.00411937400672113,0.000669320244786942,-0.0034678594687233,-0.00122355769831817,0.00327923700935173,-0.000592638145727076
"2777",0.00651910764905361,0.0133359767097359,0.00316159169770835,0.00958394549874164,0.00168926912849909,-0.000668872554844935,-0.00811931688988754,0.0071044170839496,0.012117322829762,0.00652416725529137
"2778",-0.00341840751220879,-0.000809832552305823,0,-0.00383744260310526,0.00417607779363371,0.000478164602889963,0.00272858865320691,0.00316229281422697,0.0016540564087435,-0.00471419813690632
"2779",0.00953168674713378,0.00445794798908183,0.00803665921042351,0.0131791905986414,-0.00135959504084604,-0.00219843583229606,0.00712702927731268,0.00703217431553438,-0.00809938677517319,0.00118411653188644
"2780",-0.00168080053869735,0.00100867924358861,-0.00844146655279188,0.00120061520482584,-0.0092896982864964,-0.00316117751315892,-0.00977850132881963,-0.00120419558595786,-0.00221973998905778,0
"2781",0.00454961500703988,0.00483683741280316,0.00630613761349541,0.00819503813308597,-0.00525423797159696,-0.00259491471454931,0.00649670305940764,0.00120564742126072,0.00444936433776144,-0.00177407408737407
"2782",0.00813097113674321,0.00681907301840434,0.00422992588608606,0.00574940251877343,0.000975164321208588,-0.000385265244573385,0.00813335595282361,0.0065009862814156,0.0018193640534625,0.00236963602636964
"2783",0.00212249178964119,0.00298795529780072,0.00608426347039104,0.00473101198627068,0.00430263071509795,0.00289171368555996,0.0138299786574623,0.00406739713447579,0.00497431496290068,0.00709240651970733
"2784",-0.000388230917151677,0.00317769428254255,0.000310146823091051,0.00843642148606816,-0.00541592703044214,-0.00192211628315209,-0.0035364950641662,0.00619476902038785,0.0121778992157284,0.0105631140112774
"2785",0.000423518132113498,-0.00395941969079128,-0.00480550393537027,-0.000583770075023082,0.00820874091395485,0.00221457461147345,-0.00190130522165799,-0.00331540132791674,-0.00667547144802505,-0.00580700294982217
"2786",0.0115779025928588,0.00795057205544625,0.00732086461518611,0.013821396488829,-0.00370800950781169,-0.00297860806043682,0.000380833573938588,0.00855315826557645,0.000781480028276382,0.00759347409706135
"2787",-0.00663000117813961,-0.00986001284778293,-0.00850468114742009,-0.0151690142502826,-0.00695844889623898,-0.00250527201863604,-0.0128220136151295,-0.0150764662755291,-0.00562199547627107,-0.0028985109481735
"2788",-0.0102569153308684,-0.0067715400852375,-0.0127885394460747,-0.0136479190705624,-0.00586670832229597,-0.00231891655833294,-0.00540125331678731,-0.00478372874787403,-0.00431876724489622,-0.00697676784298473
"2789",0.000496836041106841,-0.000200402693238066,-0.00568724902696516,0.00869727454485747,0.00590132970237356,0.000290693003355269,0.0157743811054367,0.0108149952422565,0.00670346198651117,0.00117094409959151
"2790",-0.00113525755868338,0.00180507512613026,0.00492537471805199,-0.0135213467322498,-0.0144927698134225,-0.00515845344665611,-0.0166750628175851,-0.0116503414164555,0.00329028588656044,0.0099413840415421
"2791",-0.0217698798367458,-0.0248248640146986,-0.0147035225530051,-0.025625756448228,-0.00927939922867027,-0.00370385921677407,-0.0102266014873212,-0.0204472146673327,-0.0131178879376496,-0.0162129851678451
"2792",-0.0418225545453044,-0.0412646485192778,-0.0473363469251706,-0.0350662107814823,0.00944991673422257,0.00821759855046222,-0.0321736034037352,-0.0351178411389318,0.00253184589391431,-0.00941735710162106
"2793",0.0197023434401884,0.0220556884553873,0.0242547442562946,0.0325373398520228,-0.0062132474849097,-0.00436628398021977,0.00351349626525943,0.0132348734742962,-0.0104964249901067,-0.0059416896181449
"2794",-0.00542489176722516,-0.0121517686053776,-0.00888019677985896,-0.0315120224675709,-0.00950331059155485,-0.00292359076925397,-0.00390543483515582,-0.009796672721473,-0.00470566289772678,-0.0113568727483593
"2795",-0.0375089137333084,-0.0250264282474072,-0.0296997128071651,-0.0346504016659065,-0.00109381815105158,0.000879688833127501,-0.0294712079978379,-0.0228308400889325,0.00152257391199151,-0.0102780351854992
"2796",0.0150214117995702,0.00348048636594633,0.0100889805270943,0.0159773120668247,-0.00631906169971097,-0.00175805602469392,0.0207549698767009,0.00882646071074999,-0.00168031681036196,-0.0146611405460728
"2797",0.0146846660665334,0.0123564131397067,0.0194684686997029,0.0157259614243384,0.00440902403930932,-0.000293129743374476,0.00300209488930214,0.00823471055392178,0.00480889648494576,0.00619967137823907
"2798",0.00248733393719891,-0.00214140580614963,-0.0122883242708391,0.00763516238601647,0.00447405517015786,0.00166352749461329,0.00761918674191642,0.00306261206724301,0.00566322870710945,0.00184840363382421
"2799",0.0134963761854321,0.0199571101424367,0.0151311953525595,0.0250474007792596,-0.0110933839444292,-0.00605713158724075,-0.00486095297925027,0.00610710654288149,0.0170526171152821,0.0153751344041695
"2800",0.0127598882981752,0.00736380420763272,0.00480280521912535,0.0205338095279526,0.00339917338773432,0.000294821034051207,0.00990488019555813,0.00354063665251947,0.00116984328690162,0.00181718054121949
"2801",0.000292917826434147,0.00104428214044217,0.0153288605567954,-0.00321928800575311,0.0054206024646275,0.00235825337089257,0.00846446040730386,0.00579641352591764,-0.00327158423151652,0.00181375993405042
"2802",-0.00626122871828161,-0.0110577143035286,-0.00811691670498738,-0.0137262686143003,-0.00438041700682612,-0.00107829967302409,-0.0123901562364159,-0.0050113532290692,-0.0134417084514044,0.00301758450131029
"2803",-0.00497404264233003,-0.00443047604907354,-0.00998352771476296,-0.000818766045457164,-0.0122684602846409,-0.00294412522603649,-0.0165924812265242,-0.00805832965616993,-0.00459437586492994,-0.00120347674362009
"2804",0.00129619231703315,0.00508590529229291,0.00462882068819193,0.000614534655617449,0.00299835352905076,0.00137804313612877,0.00932796732293784,0.00279254138843243,0.00509310026760779,0.00903620732628263
"2805",0.0159391402531959,0.00674667593824418,0.0146452853615355,0.0178096988586951,0.00888178251289551,0.00383327996454774,0.0169883397774153,0.0151899645217324,-0.001266856660328,0.00656719708467035
"2806",0.0116123543712321,0.00649223009999766,0.0129745075444161,0.00925184583840655,0.000338778181010246,0.00117493448386674,0.00347431118028307,0.0107230530321545,0.00245757097239219,0.00533812706251435
"2807",-0.0124865370665703,-0.0158136912574516,-0.0136087683606799,-0.0290953901846861,-0.00143870289538772,-0.00312968285326709,-0.0210412262005419,-0.0217121296185998,-0.0104389089072101,-0.0100296031652974
"2808",-0.0101300138997269,-0.0109935916610695,-0.00876475423862078,-0.0143677679064963,0.00635587092189849,0.00235448004158445,-0.00244850152606946,-0.0103405938342794,-0.00103889557353709,-0.0107270933030973
"2809",-0.0145409669801539,-0.0106883546840206,-0.0289832054392388,-0.00187414263185781,0.00682631703694137,0.00430355815861128,-0.00313676978322219,-0.00305804617034944,-0.00223999200000002,0.00180720426467462
"2810",0.00515511781751465,0.00108038528617782,0.0112984599482904,0.00417273741213275,-0.00812940749703039,-0.0037091872968904,-0.00177836997715441,0.00996911411950108,0.00537201727572145,0
"2811",0.0115579873326033,0.00669112296369434,0.0045023086523146,0.0014544198935158,-0.00270372784900563,-0.00127362845820178,0.0112375006508145,0.00202482400049386,-0.00167476674116562,0.00601333289763395
"2812",0.00253498226392446,0.00578909015645723,0.00614202784132534,0.00933608881385672,0.000931836298877498,-0.0000980033750980214,0.00636952138332614,0.000252693053084174,0.0107844623741811,0.00358632258656688
"2813",-0.000366350414416905,0.00255800625581015,-0.00841435346047192,0.00102774565307184,-0.00110027382820854,0,0.00511722047326901,0.0050506706706932,-0.00640162812298772,-0.0107207044128849
"2814",0.00483887436863584,0.00170119017867298,0.00615640422717045,0.000205320823285948,0.00576222239020363,0.00206012692204616,0.00509083890269513,0.00427135479059726,-0.00238627901379029,-0.00602051145286409
"2815",0.0174025037131,0.00466991529880945,0.00248042124046899,0.0213507954181713,-0.00657160824602898,-0.00215386658265126,0.00626531741245917,0.00150082436755539,0.000956809136609893,0.00969115162118062
"2816",-0.00125508131415064,0.00169013696587705,0.000989857290128127,0.00241210281654824,0.00576690370556943,0.00235487856923511,0.0050335169497433,-0.00299758078448242,0,-0.001799615516479
"2817",-0.00646270448860498,-0.00864787870793438,-0.00164793134925645,-0.00902342991242167,0.00505960313443699,0.00166392085975708,0.00158162042007581,-0.00375859403737833,0.00191172533127504,-0.00300482847068939
"2818",-0.00513170219308723,0.00255319852837865,0.00429177951753479,0.00161872113413786,0.00880945635310715,0.00195459748911131,0.000789779163861137,0.00653921373956834,-0.000636047071363111,0
"2819",-0.00108973725557948,0,0.00197240228831741,-0.00363621525787683,0,-0.000390002086896102,-0.000263005179406806,-0.000749360093130869,-0.00636431996096221,-0.000602764527766642
"2820",0.00108458684342039,0.00190985836480961,-0.0044292073220864,-0.00223047805664389,-0.00357640955476557,-0.0011709314340691,0.00591888548235242,-0.00248824591425423,-0.00240195352438821,0.00361883050760348
"2821",-0.0135304993287068,-0.00635445773959964,-0.0169714525681043,-0.0107700805210251,-0.00317155454556406,-0.000976957504694842,-0.00928362277619488,0.00428307978547204,0.00216697435259983,-0.0066105484132043
"2822",0.0017007842083554,-0.00127908258954035,0.00569905548109495,0.0110929159903432,-0.00401895649234985,-0.00195566239455869,-0.000791860821507395,-0.000501503334919939,-0.00448470398451106,0.00665453856253961
"2823",-0.00191920687815272,0,0.00133330351270611,0.00589173898113371,0.00109271936001853,0.000685794430111741,-0.00766097932729981,0.00175708865813551,0.0174563996051227,0.0180288471202825
"2824",-0.0249973209387773,-0.0217715705593039,-0.00915454321140441,-0.0333265085420358,0.0099094571566205,0.00411201819745366,-0.00579769030153066,-0.0122778466169848,-0.00395319408713168,-0.00767416064361603
"2825",-0.0213145041508098,-0.0065459836358891,-0.0209977126262528,-0.0202675164362683,-0.000748638389691969,0.00136502564273511,-0.0159286877586873,-0.00659564567232429,0.0129385454928113,0.00892313813065582
"2826",0.0273591649347669,0.0197672540760314,0.0142415608252715,0.0324163483180913,-0.00382770238329122,-0.00272603490075485,0.0126198615049742,0.0114915072653132,0.0052503565139852,0.00058967534721921
"2827",-0.0170118362612847,-0.0105535830757678,0.00236843462170078,-0.0181781207626273,0.0106925265587303,0.00566261162341419,0.0027094304209867,-0.00580660024893676,-0.00615841133581552,-0.00412480965262829
"2828",-0.00295493421349857,0.0065303796231162,0.0113079944740968,-0.00504944288558262,0.00264474080897648,-0.000193989597214173,0.01931908202976,0.00761801099708914,-0.013804965311867,-0.00414207687878376
"2829",0.0127778389850373,0.00843423854205994,0.0126835984613056,0.0209346046901102,0.0048637123783899,0.0020393546334081,0.000265062975328689,0.00856851907407075,0.000477197157149556,0.00891265673453767
"2830",-0.0215847886887096,-0.013939609407268,-0.0201054631628766,-0.0180198102730161,0.00197286237821626,0.0010189834186185,-0.013780225462104,-0.00849572330686788,0.0116861514294764,-0.0135452839627221
"2831",0.0128171877627909,0.00587211742066818,0.0126135913798595,0.00991353945848639,-0.00771237528531332,-0.00320032515399005,0.00658327957765459,0.00579647222828417,-0.0075436035275247,0.00537306070353027
"2832",0.0106990354267491,0.00410811772232011,0.00099644254870479,0.000417762201778915,-0.00206726128464108,-0.00058342646527354,0.0112119509356201,0.00927070807644581,0.00118760092190962,-0.00415671294288755
"2833",0.00789190284875008,0.00968994385817634,0.00497758012114691,0.00250510943547244,-0.00745727076365854,-0.00253100350414481,0.000924050094627704,-0.00099297357254069,-0.0051403243607826,0.00477048083169485
"2834",-0.0222859222121284,-0.00447859632884196,-0.0156843187168947,-0.0195750622325752,0.0109360810757486,0.0043914276168513,-0.00896736984976554,-0.00422465172060682,0.0046899521934034,-0.00712168600849572
"2835",0.00492843942366261,0.00921174620786469,0.00888969489488134,0.00106201835209885,0.00165157204514599,0.000194662002827917,-0.0017300406055123,0.00698764165533183,0.00340217583196578,0.0125522520913601
"2836",0.0159005920345698,0.0123114222438756,0.00548623707248774,0.0195203932629966,-0.00181371991278123,-0.00174872067910914,-0.00386541481472669,0.00669147507440204,0.00236558113862162,0.0171191926377148
"2837",-0.005242373276232,-0.00670987268459877,-0.00248007982592979,0.000416196649284384,0.00355135473202961,0.000973070210652072,0.00227468552165599,-0.00147709166388754,0.00778790101192817,0.00754505613080703
"2838",0.00822710578596686,0.00654422008126976,-0.00165761187242841,-0.000416023501696894,-0.0073244924966287,-0.0035970533618962,-0.00947924240354114,-0.000246593058474409,-0.0116306142250363,-0.00403226212851959
"2839",-0.00293297530142211,0.00167775277087068,0,-0.00998952921878815,0.00232142471710328,0.000878006223317351,0.00350452576046112,-0.000739736261498591,0.00655499905492807,0.000578361080894707
"2840",0.00822146922133227,0.000628281880856729,0.00282252601279298,0.0012612107313581,0.000330763711772208,-0.000487383824080645,0.00483541735810378,-0.000493531982141193,0.00141231858954072,-0.0034682796207488
"2841",0.0106985231423409,0.00732356264040845,0.0038079585382258,0.00209950994584007,0.0027284573092563,0.000585129511200266,0.0129662266939281,0.00691331079030877,0.000940241344673742,0.000580157907066337
"2842",0.000740197529742748,0.00332377432130082,0.0067623723110668,0.00859002657175023,-0.00799850715897854,-0.00389872110948553,-0.00171543437867305,0.00294284520007859,0.0007827632093933,0.0185506490623992
"2843",-0.0055473141250818,-0.0043478545601614,-0.00376803216165789,-0.00581631830006712,-0.00814628107788773,-0.0027401241096674,-0.014276383338426,-0.00537913877022222,-0.00195541653430453,-0.00398412652387103
"2844",-0.00847953486043385,-0.00270332573045351,-0.00197351159736281,-0.0125366749176077,-0.00720754637925392,-0.00333627067602515,-0.00858272171758989,-0.00147482895766837,-0.00760188883388535,-0.00171426242459438
"2845",-0.00014998081602402,-0.00125099056646294,-0.00131814502729155,-0.0080405679489719,0.000253071933434379,-0.00098470680739704,0.000676625467776582,-0.00664699686058978,-0.00797594585744166,-0.000572402055533772
"2846",-0.0134672452037315,-0.00501045235724606,-0.00362970466154733,-0.00469287042546063,-0.00455738857559507,-0.00118281289278377,0.00243302543451351,-0.00148711714873273,0.0048559145473035,-0.00515456898568611
"2847",0.00247144453217363,-0.00356701131508119,0.00314625122559131,-0.00771534359810444,-0.00669751986338518,-0.00217018394397761,-0.0021574322372081,-0.00297818188932641,-0.00649607051027323,0.00172709207715172
"2848",0.0101658922039793,0.00568540698669628,0.00610755609287872,0.0144708468842485,0.00699889903521633,0.0028674758820062,0.0121620109733678,0.0089617173225407,-0.00350851595539381,0.00517234311863457
"2849",0.000938698098005508,0.00125640766683621,-0.00278918374047554,0.00617408312813961,0.00771321700563576,0.00167618955519577,0.0129506468595189,0.00542816161635407,0.00424100980842601,-0.000571629824671294
"2850",-0.00769048591767096,-0.00460057962359028,-0.002303359303099,-0.0071941712984992,0.0017664187703903,0.00108268715137672,-0.00303151721850203,0.00147249166396879,-0.00725102788844623,0.00457659625192264
"2851",0.00177688120396402,-0.00546219613626742,-0.000824534834878099,-0.00490204690536844,-0.00360166494424841,-0.00156646460227294,0.00700687456401239,-0.0019603795068539,-0.0070631433361632,-0.00569480027258995
"2852",-0.0067174838946753,0.00042249561953267,-0.00594155324906209,-0.00792447880160541,-0.00109794196248791,0.000197460225978663,-0.00341341363338099,-0.00785661204098609,-0.000484981007881191,0
"2853",-0.00220384398124596,0.00358942628389314,0.000996128933526963,-0.00215888707950085,0.00448096268575893,0.00256453612982743,0.00039529667941185,0.00470175505652182,0.0050950019394258,0.00630014665445522
"2854",0.0129466049362443,0.00189356309769595,0.00729806023842317,0.00454354450430627,0.00151497642998355,0.0000985041952128451,0.0105345235924366,-0.00123149739599049,0.00209206631873249,0.00682990607890632
"2855",0.00338328090238793,0.000840000474134239,0.00115267907295102,-0.00581532986334188,-0.00159676868769287,-0.000491673944468918,0.00547318014666565,-0.000739736261498591,0.000240878430697755,-0.000565341543789177
"2856",0,-0.00125886498712691,0.00312496652650052,0.00563263581316242,-0.000925821585779696,-0.00167345809970088,-0.00492499643701338,0.000740283876325742,0.000160520189451674,0.00282807382389816
"2857",0.00966571849074005,0.00693271942051488,-0.00852590845900003,0.00193867226126043,-0.00598212337029713,-0.0022675476166174,0.0061214110726806,-0.00271268558521198,-0.00208679676015089,0.00902412904987493
"2858",0.00935045536739931,0.00479869110728837,0.00578796968773432,0.0208558047598593,0.00805238669152608,0.00207508294167136,0.00919098646539029,0.00642939946319099,0.0068366282178618,0.00503079018948172
"2859",0.00305120604265796,0.00145340210156064,0.00756327330858619,-0.00168479461620408,0.00252258577471354,0.0000987173324515922,-0.0041047490020697,0.00147399165264828,-0.00143792938169041,-0.00611782543922279
"2860",0.000476663507810393,0.000414787574506414,0.00554832719605325,0.00126571181804835,-0.00528395755849287,-0.00216928907521763,-0.00734157817722192,0.0031894479263963,-0.00408001599999996,0.0072746624522757
"2861",-0.00688699372627111,-0.00518148095950044,-0.0102240047666762,-0.0206489320005321,-0.0113830490730061,-0.00553461365711583,-0.0147917236779606,-0.012472543980898,-0.0161458352662196,0.00111115316920229
"2862",0.00420497134289088,-0.00083328396554061,0.00295131851360142,0.0150602791200685,-0.00383785988125485,-0.00208662130145265,-0.00289731656817793,-0.00470516381472974,-0.0015512899685346,0.00554942804543024
"2863",-0.000844637002328064,0.00291912603025479,-0.000163481542810096,-0.0152607927168661,-0.00505123934832974,-0.000597493684806882,-0.00515129886557131,-0.00497635557423293,0.000572409840768451,0.00110373765033045
"2864",-0.00249985538612685,-0.00374224746389085,-0.0024526410570852,-0.00839421655004813,0.00860496850826964,0.00388578718175236,0.00225707847802115,-0.00300086610746475,0.000408654785807094,0.000551146903571942
"2865",0.00751836097355518,0.00605174980950562,0.00114750798826813,0.00607763164531283,0.000511906490094249,0.000694901338551546,0.0107297961424841,0.00652120300004722,0.000571840517217925,0.00771362090786609
"2866",-0.0027801938404447,0.000414849193183686,-0.00229224961897145,0.00345189758070674,-0.00153493372774549,-0.000396697207029617,0.00131078646119254,-0.00249195514913447,-0.000571513702526616,0.00109347875985599
"2867",0.00275124645802882,-0.0143063732230067,-0.00393819547255392,-0.000429909619510838,0.00725942156776904,0.00456444266486056,0.00850791233352677,0.00174883479982335,0.00106198019567105,0.00546159048228656
"2868",-0.00204845089480854,-0.00294482576542765,-0.00609548206418242,-0.00537739148905436,0.00797015150838276,0.00256806566769097,-0.00246606864380683,0.00174569624879584,0.00856858977828789,-0.00651827470529265
"2869",-0.0023827112437339,-0.00886088469226887,-0.00331515498710533,0.0041090000804036,0.00622491614857767,0.00394109239747675,0.0033827837995315,-0.000995920165647313,-0.00307465824337438,-0.0147621883463144
"2870",-0.0115012311875856,-0.0266069857372813,-0.00665227735747875,-0.0232609571246974,0.0219026851803217,0.0107946055492485,0.0029823807299274,-0.00971827208121467,-0.00016230013929297,-0.0094340048311472
"2871",0.0133447766506507,0.0177126810783979,0.00703168953268207,0.00793821220651414,-0.0067081622932863,-0.00427176694133746,0.0126698296061372,0.010317092536493,0.00146116565531007,0.0128852670219088
"2872",-0.00612589927700047,-0.00429742089527396,-0.00681633633891265,-0.000437502734392026,-0.00164727350150851,-0.000487334428396768,-0.0017874637144446,-0.00423420707002842,-0.00218857901786706,-0.00276550571138057
"2873",0.00981782294851441,0.00820034690831828,0.0068631176571976,0.0140075959969066,-0.00528357378702704,-0.00369486504646666,0.00345313030416206,-0.000250056149049493,-0.00495532095784434,-0.00665559702864238
"2874",0.00475148838461092,0.00256831771394261,0.00598496395432369,0.0101443832648258,-0.00723197444420209,-0.00353189404291365,0.00879422800768648,0.00850635067395289,-0.000979631006280179,-0.011725247698573
"2875",0.000727402407743272,-0.00170799988958792,-0.00181782583998613,-0.00769219656948505,0.00234457202902827,0.00255974954842508,-0.00126338751093302,-0.000992262888789841,0.00392248907601966,0.00169489199511852
"2876",0.00836062615054889,0.0100514597660437,0.00430462116181451,0.015073160601941,-0.00810307445040603,-0.00402608041583241,0.00113848978881514,0.00645620004679714,0.000569800579077073,0.00338416449252255
"2877",-0.000108194146018148,-0.00804575239772232,0,-0.0152735652070265,0.009685106005622,0.00423984326536275,0.000631773571260652,-0.00764849388090894,-0.000488097957827893,0.00393474064972654
"2878",0.00295639628112343,0.00128072073713725,0.00296732272794431,-0.00193874021252616,-0.00300279045189233,-0.00137472382429826,0.00290442248514755,0.00198902336101203,0.00122090996890023,-0.000560017988806005
"2879",0.00133015897087052,0.0100191359509798,0.00312298023295465,0,-0.00184053780009286,-0.000983225879385707,0.000251813154692471,-0.00198507500046274,0.00178848058225367,-0.000560216466350849
"2880",0.00129225472264971,-0.00654283923743459,-0.00622639623611476,-0.0025902503771017,0.00025140308641447,-0.000590497741857265,0.00503519512299011,-0.0044754303805894,-0.00332713616829172,-0.000560415101785283
"2881",-0.00319104784308588,0.00212448257383535,0.000824347530323344,-0.00670846337066688,-0.000502539911727662,-0.00118170349725233,-0.0201652261411923,-0.00174816954485557,0.00301255495847585,0.00392579808687055
"2882",0.00251792099557147,-0.000635982325706164,-0.000988484255802557,-0.0067538624227701,0.0082995240746282,0.00315506380066299,0.00997060166110142,-0.00375272358849077,0.00154229236882375,-0.0111730327424138
"2883",-0.0012758392254244,-0.00615188463356386,-0.00527704688541009,-0.00789651522607793,0.000914572025654925,0.000785991741264036,0.00101239902725325,-0.000785802401078062,-0.0165342928319248,-0.0242939171124082
"2884",-0.00205666977649288,-0.0091783205456758,-0.00729431003484171,-0.0121600295916819,-0.000913736347952332,0.000491186644683728,-0.000885036886331014,-0.00532586615848807,-0.00189545910319633,0.00868564270287542
"2885",-0.00383292351352926,-0.00844301625929922,-0.0106025435886629,-0.0110384897774766,0.00582029323787103,0.00265018218925905,-0.000126450138779655,-0.00535441175078244,-0.0025596399755623,-0.0103329868542164
"2886",0.00170595555927333,-0.000222243720307547,0.000340194235066926,0.00432798546286106,-0.00876239731692996,-0.00323063473737917,0.00974562365617193,0.00281980400673132,-0.00447020684262733,-0.00116019641551013
"2887",-0.00626880974665001,-0.00778289768124085,-0.00374096895489739,-0.0140620047128914,0.00525390002703752,0.00265174410450619,0.00513918072593555,-0.00460126063822308,-0.0017462081864924,-0.0075492592332711
"2888",0.00182320704859218,0.0136708385401572,0.00494971684439172,0.0103518570197556,-0.00008307863631829,0.000195957988088358,0.0063597087888283,0.00950183513247316,0.00241560177220479,0.0198948260359761
"2889",-0.0136127947074606,-0.0148129732975072,-0.013586917624913,-0.0134334187857085,0.00224027976021124,0.00137106087349181,-0.00346944129962279,-0.00661411584684679,-0.00373938021403952,-0.0114746066791805
"2890",0.00221414466386416,-0.000224431859121799,0.00585385834586627,-0.00392351231522559,0.00140716355501413,0.00048909789647289,0.00395499002474908,0.0040973766132455,-0.00525479193639833,0.00986655672432346
"2891",-0.00828440803937569,-0.00965215228217298,-0.00667574159840878,-0.0192307631799801,0.00942398258096588,0.00381217890122509,-0.00537782668705877,-0.0119867610149303,-0.00570182784333684,0.00517234311863457
"2892",0.00571740815070676,0.00249325309116055,0.00120622953537253,0.0085046360443537,0.000245698158901853,-0.000973842709021011,0.0106878767264156,0.00309752795965013,-0.0030359334957677,-0.000571629824671294
"2893",0.00143981564996354,0.0108522814175827,-0.00327012986893371,0.014991901655999,-0.00343894637090714,-0.000779556241574997,0.00248821168137048,0.00720525649684145,0.00363729484319664,0.011441608389076
"2894",0.00213808323992204,-0.00715719027888451,-0.0158867186716306,-0.00992399385231391,-0.000782238804042157,-0.000684329342301893,-0.00595680796995435,-0.00715371216578231,-0.0100295236404632,-0.020927723011414
"2895",-0.00353133354905932,0.00585717731587532,-0.0012283139585213,0.000699351833970407,0.0053563402499972,0.00254287927503771,0.0074904273138201,0.0059187679448971,0.0101311340893167,-0.00115526692314427
"2896",0.00815794282177107,0.0132139276411276,-0.00158119526929035,-0.00256244119364391,0.00286887920832712,0.0000975180316087343,0.0130112818838837,0.00690710056750121,0.0033712683797511,0.00578367033561245
"2897",0.00845821365034061,0.00486280262766225,0.00651069783435787,0.0137786815979142,0.00326923400573786,0.000877839585639251,0.00415882895289665,0.00685971979302602,-0.00159598484008439,0.00460028213185626
"2898",0.00900442316554084,0.0063793741323166,0.0138111934818705,0.0179682246578181,-0.00643557672148698,-0.00253395770930565,-0.0088925665005517,0.00454207545283847,0.00243985358876109,0.00515173632649257
"2899",0.00359827498500942,0.00240433131790208,-0.00379381451787619,-0.00226293964438407,-0.0000821904326460121,-0.000781556375471837,0.00307294932642144,-0.00276325233844732,-0.00184642884017738,-0.00227787321992068
"2900",-0.00731426846984984,-0.0183165532169245,-0.013847978993315,-0.0195055058245853,0.00385419364353234,0.00205328265603799,-0.00306353523787573,-0.0130981687954941,-0.0108467249642648,-0.0348174624831071
"2901",0.00906585185982434,0.00888485406674011,0.00105316887974105,0.0136479036866912,-0.0000818050681147264,-0.000390014440821096,0.00294995351443905,0.00535973372072895,0.00416523294938154,0.00532240485517366
"2902",0.000787572131371927,0.00286218790593917,0.00929340896055453,0.000684573568380253,0.00253257575075949,0.001659323684291,-0.00343124770261916,0.000507855448876438,-0.00440189632782273,0.00176480282097224
"2903",-0.000894157917387783,0.000439016598250186,0.000347481730034183,-0.00547312785178355,-0.00415587067523981,-0.00165657489034077,-0.00455010408596646,-0.000507597662637638,-0.00051014369092639,-0.0211392979429703
"2904",0.0040452566923137,-0.00175534146653578,0.0088571343194126,0.00733779152586345,-0.00188208362391251,-0.000585862097964185,-0.00531186349338608,0.000253927724438219,-0.0108039469807585,0.00119974367765274
"2905",0.00210365010658675,0.00241798164218276,-0.00154927736587518,-0.00113822576932954,-0.0040169425722919,-0.000781337388150338,-0.00471940844695029,-0.000761244978765729,0.000257989338303899,0.00898741846514817
"2906",-0.00377155534964879,-0.00350882950969988,0.000172387353531755,-0.0123063082622605,0.00633797194117847,0.00273699149089568,0.0101073391753534,-0.00558803879961378,-0.00429885657809059,-0.00118763226939633
"2907",-0.00114285056650021,0.00572192521330295,0.00310298746917725,0.0143055166666228,-0.0122689554289368,-0.00350955713239554,-0.00840018242834151,0.0109834255019154,0.00647612479882786,0.00713438888152895
"2908",0.00185919030386028,-0.00262579524367568,0.00498359939304716,-0.00659697637731194,-0.012338621131966,-0.00489113463822133,-0.00249172598794001,-0.00480063599645797,-0.00480437551139967,0.00354192497063477
"2909",0.00503213528995383,0.00680105438023548,0.00410402422008316,0.0146553970809096,0.00343776324625766,0.000687897111421032,-0.00487060872552214,0.00330057181879351,0.000344836206896515,0.00529404521019172
"2910",0.0085224473504828,0.00740909862630712,0.00647136094667911,0.0162490921267611,-0.00158760196966401,-0.000687424234276035,0.00815768472681722,0.00607278466897876,0.00551533087284284,0.0134581601662647
"2911",-0.00235896966808713,-0.00605654763412311,0.00253808233543062,-0.0111037245934639,-0.00192499584386296,-0.00108168139520237,0.00273872331094394,-0.00829984049347332,-0.00779913438464175,0
"2912",-0.00677628258184326,0.00195858074650701,0.00303797771750203,0.00359309604217528,0.00167704379193734,0.00157458827869195,-0.00968357077244886,0.00152167604528208,0.000518312184114356,-0.00404145601756001
"2913",-0.00522344962191823,0.00260640409212165,-0.00757198419526428,-0.00156630471810926,-0.00343203396400982,-0.00127728885288769,0.00137886984486824,0.00177284942456502,-0.001554001527169,0.0057971412257396
"2914",0.00492911523773065,0.00411597121832408,-0.00762968680031517,0.0053788429181918,0.00545995354050399,0.0013772649664312,0.0171508806615657,0.0045498825977528,0.002939870247473,-0.00576372808007275
"2915",-0.0016704935896461,-0.00755106247583337,0.00649235099316736,-0.00891672968623669,-0.00814688713309564,-0.00236254608323949,0.00332304683649753,-0.00603930862187485,-0.00732820945474966,-0.0144927933996526
"2916",0.00544764042257273,-0.0091304033433266,-0.0056016578773358,-0.0132703313464081,0.00143514471901884,0.00118422869328816,-0.00331204076989478,-0.00278493882566933,-0.00538476641814112,0.00588239354001052
"2917",0.00428483338734642,0.00197445693757392,-0.000170750808167863,0.00775026933724754,0.00497346531663689,0.00256246591868936,0.01181528481015,0.0040620100987645,0.00349284850225762,0.00350872377936784
"2918",0.00366709653712971,-0.00459826872031011,-0.00751231566041777,-0.00769066461509815,0.000587199377668712,0.00049178447865339,-0.000608161420662112,-0.00455103430698256,-0.00513397154775463,0.00174822784108608
"2919",0.00330235584121263,0.00791915753652983,0.00842932844193856,0.0102575434371421,-0.00519732793782435,-0.00206365614261672,-0.00352955675325184,0.00330190267591113,0.00227406625952842,0.00756249299486456
"2920",-0.000420155899479635,-0.00174585481003298,-0.00102352492264934,-0.00135379536807212,0.00101109646797903,0.000886413053182933,-0.00598519070033554,-0.000759518348429911,0.00279263470783264,-0.0121246057469363
"2921",-0.00136610318108255,-0.00349808934594753,-0.00375686944404663,-0.00293705805499078,0.00841806558688529,0.00275436217343694,0.00122881828111576,-0.0035468357891929,-0.00147947083876176,-0.00409111864171874
"2922",-0.00670011352552313,-0.0223782137557023,-0.0143983515651468,-0.0213008219146434,0.00726280476213281,0.00431667578330952,-0.00895913882732635,-0.0142386484245306,-0.000435732969073177,0
"2923",-0.00374347179290946,-0.00269313559661877,-0.00591303161338774,-0.0164388788545115,-0.00207205116752596,-0.000293136468350497,-0.000495426996524051,-0.00464282835928109,-0.0150841657496876,-0.00528167780563416
"2924",0.00638062001702244,-0.00180009255852376,0.00402373390710764,0.00612054807698414,-0.00224220296704625,-0.000977074488745511,0.00545155381040474,-0.0025911848434359,0.000973804895306296,0.00176976566726261
"2925",-0.00746731681526347,-0.0171326916457107,-0.0121972061268161,-0.0287787587415663,0.00582650890192649,0.002445262435951,0.0075170300777978,-0.00545605119394166,-0.0166268506235074,-0.0217903474683254
"2926",0.00809148259901393,0.0071102927387634,0.00546835125206191,0.00626354753842007,-0.0000827585882041681,-0.000292793246562728,0.00807235191480382,0.00705325461426698,-0.000809461267929579,0.00782656574689478
"2927",0.00352035273774032,0.00592110946999935,0.00333332767644468,0.0105339126053279,0.0012414471810156,0.00039055581693459,0.00897847547096542,0.00648505059646309,0.00927091825870252,0.00418166710267975
"2928",0.00213987506005053,0.00701834738735463,0.00402169519788687,0.00450134324093443,0.00669537044528035,0.00312184401423887,0.00156315088339798,0.00670117138905835,0.00499424788176883,0.00178462762613107
"2929",0.00234526164362037,0.0107913801206971,-0.000174200325966156,0.0127357691723415,-0.00336660901412522,-0.00136154046911463,-0.00672332726549529,0.0017921341737861,0.00292834319055202,0.00178144840409455
"2930",-0.000593722792776363,0.00333624944292832,0.00418051452505774,0.00791805269647239,0.00395460301806838,0.00185035156065072,-0.00556046321258208,0.00178884137823965,0.00221199793519733,0.0142265489565536
"2931",-0.00132769118155462,-0.00753720921266809,-0.00416311058080521,-0.0161735909090701,0.0015592346226696,-0.000096905359134869,-0.00218807231230755,-0.00612259008104488,-0.00944645562231283,-0.00175333656073662
"2932",0.0060182295122424,0.00826451794918714,0.00348373521676471,0.0185532006761251,0.00196631905972411,0.000291357763889888,0.00511657855547032,0.0048770042399584,0.0174688685597737,0.00761113664734459
"2933",0.00789547024400949,0.0132921532078663,0.0151015335874842,0.0142956204977316,-0.00572394498938111,-0.00223550869315225,-0.00181802824082833,0.00791822095932027,0.00376657309857831,0.00348629761126173
"2934",0.000483022170055136,-0.00174918119620882,-0.00307792578083277,-0.00363720253512789,-0.00600390627219072,-0.00224020499702215,0.0106847647547677,0.00126692710029341,-0.00794132150942739,-0.00405309730294123
"2935",0.00538078742641335,0.00459918468149234,0.00360207070524399,0.00616004211989729,0.00132376358457265,-0.000292964734739942,-0.000960924543257469,0.00556835410252932,0.00457421710063333,0.0110464194354272
"2936",-0.00404826991507434,-0.00981027971412185,-0.00700745274503134,-0.0260770231136993,0.00214859173113702,0.00185542130454652,-0.00348730239669393,-0.0113263656805797,-0.00490366037400147,-0.00172510579944607
"2937",0.000034418000024683,-0.0112285921364474,0.00206551297911783,0.00512225272299816,-0.00230877338253221,0.000194954821718385,0.00374083840192241,-0.00152757322853347,-0.00114393700408255,0.0011520579548232
"2938",-0.00172228411634034,-0.00823866165796805,-0.0123669316059342,-0.0194579991046908,-0.0057815605244852,-0.00228507282355805,-0.0105796207845879,-0.0114737642079799,-0.00510969949590867,-0.00575372044135014
"2939",-0.00269141306836218,-0.00583745204379282,-0.010608661732083,-0.0144105592641929,-0.00266622250203075,-0.000097676567903604,0.00461733660601316,-0.004384956718679,0.00345346674931357,-0.00405098955429095
"2940",-0.00301000601739754,-0.0049683942490315,0.00228510482726429,0.000958776059713395,0.0036756520643122,0.00205543055082047,0.00387046719120687,-0.00103602950695569,0.00194141369572898,-0.00581049601876982
"2941",-0.00194338299339725,-0.00817059828053601,-0.00613823028804095,-0.00502877788020129,-0.00848925358770092,-0.0044933904097213,-0.0121687281422909,-0.00674276127906348,-0.00273029766839628,0.00233778208098223
"2942",0.00173850918334262,0.00892447655316331,0.00229397598097636,-0.00986761331554453,0.00369328559556514,0.000588658791623287,0.00634219934200542,0.00104438086618108,-0.000706535351765347,0.00349849440394534
"2943",0.00329726544369224,0.000453577826141416,0.00211269635556022,0.0021877102578749,-0.00761047636664702,-0.00362847199915606,-0.00206050232176469,0.00365148992635711,0.000618638963877371,0.00987802264203652
"2944",0.000242395342547441,0.00385398211431975,0.00193252981082548,0.00509324388332266,0.00235964304350778,0.00118100130769938,0.000850265118908844,0.00545735171705508,0.00839071711366635,0.00690439346752192
"2945",0.00591446235494697,0.00722678732238702,0.00771524546000113,0.0135136368270001,0.0015134208568095,-0.0000984233267161683,0.00594587069432628,0.00361857490445661,-0.00359110105266014,-0.0108571717928199
"2946",0.000171879046668044,-0.00224218924851982,0.0113101975962075,-0.000952384197535516,-0.00478523552141719,-0.0018677403177294,-0.00808215751557928,-0.00309046509343591,-0.00650496648198018,-0.00635450319835917
"2947",-0.00529433390747569,0.00269669693858243,0.00051623595361372,-0.0090562500343867,0,0.000196766598396181,0.00352675636901933,0.00258338601998398,0.00522035051903247,-0.00116289437072703
"2948",0.00542632315598679,0.00515457196554658,0.0239036946898419,0.00962001736592022,-0.0104597726340337,-0.00413597305393254,-0.00351436207020528,0.00669923956540996,-0.00149633833732643,0.00931320734642194
"2949",0.00106564785300312,0.00222969106137638,0.00352703553878886,0.0138161251222619,-0.00596700429874042,-0.00168139854132043,-0.0132553934231512,-0.00358317730448443,0.00387865825319711,0.0063436269774495
"2950",0.00810376366278986,0.0180199821257478,0.00267782696580698,0.0110431968543943,0.00463070689730394,0.000099010411342082,0.00998277189087737,0.00796285136842489,0.00342465762446409,0
"2951",-0.000913727558023658,0.00043702463620332,0.00216991514095666,0.00464793596539637,-0.00042661915260167,0.00039626832026407,-0.000487980555292644,-0.00789994527835469,-0.00682592999455489,0.00229223237918608
"2952",-0.00332190671311938,-0.00480551203005752,-0.00449698083657923,-0.0113346873852362,-0.0025618428793186,-0.00108912733418065,-0.0175803569225021,-0.00363363491388358,-0.000176200549408811,0.0148657296621684
"2953",-0.000927930029337665,0.00570676254228153,0.00752891112892518,0.00397740537521996,-0.00102754834331598,-0.00099098969845135,-0.0016156003462896,0.000520837832959753,0.00158633117488027,0.00225360625707682
"2954",-0.00299205435955541,-0.00152768542268467,0.00481553512866739,0.00209744488717556,0.0070277561773362,0.00327416867826469,-0.00915059433139487,0.00364501709147813,-0.00527935758417319,-0.00449707787132436
"2955",0.00279419671709302,-0.0028416106876884,-0.00264417689167384,0.00488368930950589,0.000680927776752549,0,0.00266408314408251,-0.00181584599868023,-0.00884564328582993,0.0045173929391471
"2956",0.000103292465039706,-0.0120560973157002,-0.00198836900983113,-0.00671145709727794,-0.00263651981781476,0.000494025685088051,0.0123985406369411,-0.00597721314155264,0.00633644784462883,0.0101179045278676
"2957",0.00347412438632522,-0.000443784543227688,0.00680727158259242,0.000233114132708545,-0.00734124497211752,-0.00253530280262826,-0.0082476868724517,-0.00261430698059961,-0.0016850123858636,0.018920451388869
"2958",-0.000582803990135106,-0.00532729375464069,-0.00230876034615191,-0.0125786351757077,0.00611261772587035,0.00258170915812772,-0.00138608322308387,-0.00996072915960844,0.0115483965532557,0.0032769655314917
"2959",0.000548818110525096,0.00379361414247392,-0.00876031430284863,-0.00825661886464868,-0.0173712202287843,-0.0074280137650079,-0.00694011419176022,-0.00529518033098042,-0.00395191875071776,0.00925425988695894
"2960",-0.00781572187205082,-0.0131168220587201,-0.0135066901799198,-0.0249761987618015,-0.00705397286599629,-0.00259410564953788,-0.0100380909625135,-0.0188979970428516,0.000529051323030272,-0.0107876155675189
"2961",-0.00559710487549725,-0.00698356388127841,0.000169007203053573,-0.00365949250137498,-0.00859488227069238,-0.00240101610542276,-0.00128366170294647,-0.00189907059746985,0.00281988008054612,-0.00218110757682066
"2962",0,-0.00930131679799473,0.00439412303544495,0.00146915296724637,-0.00336163208218676,0.000401099756657919,0.0132374512215165,0.00462073856346801,-0.0110720735218258,-0.00273220340393854
"2963",-0.00145920392672028,-0.00114495769254785,-0.00572107396498189,-0.00366754538905723,0.0101189123068077,0.00190458132463212,0.00215623711673119,0.00865810301825354,0.000533117109177805,0.00712324725195068
"2964",-0.0316631593085488,-0.0194863534993317,-0.0245387517141701,-0.0296931507380268,-0.0027241930539893,0.000500130761798223,-0.0150612631806833,-0.0179719806688364,0.00248666967116651,-0.0195864096426023
"2965",-0.0220264321236416,-0.0126258055047875,-0.0180430430716371,-0.0101163459436877,0.0121598848289721,0.00410001134842153,-0.0272424821594417,-0.00409741789555229,0.0256910176920009,-0.0149833186461571
"2966",0.0138883274470145,0.00189456695698653,0.00229674022630433,0.029381700311466,-0.00348211194593195,-0.00119501002887967,-0.00198145217677403,-0.00191990522817009,-0.00475035416091174,0.00788721601174891
"2967",-0.00561705818107028,0.00165442067713695,-0.00299660863246398,-0.0106726859329337,-0.000437017537151196,0.000598225030130628,0.00542685217588623,-0.00109917266765425,0.00668226138985695,0.00223597067338011
"2968",0.0218657750337623,0.01604517349859,0.0185643480590378,0.0250879471836001,0.00227250329038386,-0.0000998019998144084,0.0217219291421529,0.0198073107446226,-0.0017241120689655,0.00446184972113572
"2969",0.00017847054166964,-0.00952154904876357,-0.000694288889770078,-0.0122370241891204,-0.00592955446775034,-0.00288980272740913,-0.00489626465531778,0.00161863574435928,-0.0000863730547572272,-0.0088840601011867
"2970",-0.0144411933220425,-0.0164126865136246,-0.0180649823128983,-0.0262635890306195,-0.000350997390069163,0.00179904162337019,-0.00116532129764024,-0.00430906476739323,0.00112269625077555,-0.0112045023045214
"2971",-0.000542596351723712,0.00786647578168509,0.0021227870212448,0.00941473739094789,-0.00219368730907432,-0.00119715585662672,0.00764854476154198,0.00405727655269716,0.000776432035480168,0.00566582033804575
"2972",-0.00448872240494458,-0.00591292319831371,-0.00617832109645589,0.0108393836521843,-0.00131926068584964,0.000199454641462982,-0.0131225574474467,-0.00484933559948786,-0.00258600978215662,0.00112674514453537
"2973",-0.00509069212788504,-0.00713775220408586,-0.0115452409161565,-0.0109724766302115,0.00317019698679588,0.00259658140826136,0.00638777177902661,-0.00378982534887617,0.00587676091847511,-0.0219470914597191
"2974",-0.0302985233213612,-0.0282769595835076,-0.0319856924745601,-0.0322743888021586,0.00754916627360935,0.00537901196128798,0.0072539104703,-0.0138588153170957,0.00231982990222379,-0.00690445268593698
"2975",0.0179403243372234,0.0128235763053226,0.0148506007417497,0.0192808060151362,-0.00418172456850208,-0.00237794144853232,0.0123456077983588,0.00909367359125857,-0.0022287158502069,0.00405556430793319
"2976",-0.0175873134693278,-0.00413917782058759,-0.0128040537354562,-0.0115030546247896,0.00603651490263823,0.0044693049680391,-0.0235008495145855,0.00191142481283357,0.00317865114813309,0.0075013995081854
"2977",-0.00554035290854493,0.000244439161749099,-0.00926439600485041,-0.0173260453693882,-0.00226090581534166,-0.0000987881424155956,0.0115778872366681,-0.00327067766530698,-0.003939359525718,-0.0103091969184586
"2978",0.0148186053956292,0.00855536600843476,0.0157097395019186,0.0194738066409266,-0.00496827464633132,-0.00217548966984227,0.015046349289517,0.00464865920182511,-0.00438479072108655,-0.0052083811063095
"2979",0.0106808231205724,0.00799812935216959,0.00975869724266243,0.0108413280188648,-0.00508056308918292,-0.00247742581907784,-0.0103889051955918,-0.00816559681264017,-0.00561313456960799,-0.0133799887343048
"2980",0.0106417997542847,0.0158692085988228,-0.00237052556661188,0.035750918647101,0.000926723544785846,0.000856155488343058,0.00371274270241773,0.0148189333091115,0.0128527570498871,-0.00707537594761776
"2981",-0.00592298047950413,0,0.00566631192418332,0.00641017501899466,-0.0124328174235866,-0.00557035993941501,-0.00854593570061002,-0.00459699805888514,0.000171525340946443,-0.00237526453879289
"2982",0.0055169923331444,0.000709935293166764,-0.00363513885639388,0.002694817962686,0.0039286547485291,0.000599942268386666,0.0146660215752101,-0.00135848679383055,-0.00240033429232178,-0.000595229963322619
"2983",0.00632794289678107,0.00165559486421696,0.0113097718436566,-0.00171019175157183,-0.000622525702074772,-0.00109965952357172,0.00431092606047168,0.00788920414669092,-0.00283579953160262,-0.00416921391002356
"2984",0.0214088304093247,0.0129870921385065,0.0104617527745046,0.0188447201796276,0.00133477132687809,0,0.012624657269928,0.015654631381923,-0.0000861944149759264,-0.00239218884047798
"2985",-0.00181500492380027,-0.0114219413258506,-0.00642622794948,-0.0259428944320121,-0.0000888349689861512,-0.00140090909581092,0.00037390965239914,-0.0087698460104072,-0.00215461520429727,-0.00599530645430091
"2986",-0.00976813699014956,-0.00377258541306236,-0.0100611321817843,-0.018495646572353,0.0074659268143682,0.0039083281460317,0.00137107622968768,-0.00482560418882905,-0.0112281569461752,-0.0108564294470516
"2987",-0.0186851487975579,-0.0201182901969638,-0.0136115641135693,-0.0140702958894899,0.00652846377589866,0.00299514965971759,-0.00112017498124084,-0.00592677120494634,-0.00716281427770404,-0.00243899102184708
"2988",-0.00187120557279885,0.00748773044522344,-0.0036798753979963,0.0114678760482385,-0.000613658254639327,0.000796211635170962,0.000872205565065176,0.00785902819589124,0.000351865199652801,-0.0275061756106754
"2989",-0.00683655083627943,0.00119876057708068,0.00350882300752553,0.00604685771899161,0.000614035062323826,0.00208840168684876,-0.00174278756747781,0.00349572289369338,0.00826738808093386,0.00879950644204519
"2990",0.010436596887323,0,0.00588883474402446,0.0222890042466346,-0.000438171035292423,0.000695043658619277,-0.00623513367673567,-0.00535911814033729,0.00113396721156644,-0.00186913334812067
"2991",0.00260061734762296,0.00023950493010072,0.000731759623402439,0.00195983038653758,0.00578752921075232,0.00307426943923939,0.0120465185927909,0.0037713264725272,0.00740616905304958,0.0062422403245177
"2992",-0.0169146021047345,-0.00766095219158702,-0.00438755420008141,-0.0134475046697691,0.00278980479613411,0.00148313555820589,0,-0.00214689530917278,0.000432407876689078,0
"2993",-0.0185062207176934,-0.0176115548962528,-0.0183621001177368,-0.021561232983661,0.000347589513761459,-0.00019764193710381,-0.0106633727389087,-0.0134480498269419,0,-0.0303970519984572
"2994",0.00340764954604489,0.0135068288006506,0.0153385477487715,0.0184902527711024,-0.000347468737272094,-0.00019728505629657,0.00137871765620434,0.0111777340481065,0.00164262992379394,0.00831735623043794
"2995",-0.00667862047395595,-0.0079960903452243,-0.00368454527516271,-0.0116884161771456,0.00104325283660511,0.000592591386076924,-0.00337923073571367,0.00242650819272039,-0.000776834103427881,-0.0291878088056222
"2996",0.0161441786425613,0.01587691143772,0.0134984481807219,0.012330029070281,-0.00225809264765675,-0.00078975200889797,0.00351622866745571,0.00968256814969726,-0.00112289888026862,0.0045751006142738
"2997",0.00336447316669575,-0.00456834294192809,-0.000912233854500899,0.00695990010606296,0.0011316060747284,0.000987972801771209,0.00312849078969757,-0.000798961350244598,-0.00596681084371165,-0.00390365519694513
"2998",0.0230253347231717,0.0132848760520181,0.0131482406311618,0.0239446858383787,-0.00486918781167345,-0.0000986957088623397,0.0088574523375835,0.013063103833618,0.00374075694843223,-0.00326592898342237
"2999",-0.00218510740265832,-0.00452923865944366,-0.00342450355604973,-0.00867881125388648,0.00393189205358202,0.00256592566680958,0.00136009951243676,-0.0115789507826256,0.00312013355313234,0.00655312555937493
"3000",0.00609547239196551,-0.00574707157870258,0.000904258352552256,-0.000972664391154954,0.00374236842228126,0.00196907680377278,0.00987891433477239,-0.0106496602717474,-0.00172798516896466,-0.00455729637804392
"3001",0.0132411954982041,0.0108381903701067,0.0135525508942627,0.0202044705972819,0.00710041714814347,0.00218577803068865,0.00464660176348231,0.00188364859143975,0.00752988568868029,0.0228908020595362
"3002",-0.0324022554893663,-0.0228735085321919,-0.0369049108196652,-0.0212360533224223,0.016741335457874,0.00461733993365532,-0.0154576274853468,-0.0104752996298474,0.00609912357704245,0.000639377437478439
"3003",-0.00151715361828597,-0.0141429209945474,-0.00148099154787262,-0.00926380561669682,0.00314061850468716,0.00254233103887636,0.0250958598325626,0.0114004268225494,0.00017073086994368,-0.00830666140199077
"3004",-0.0232358117026542,-0.00964629347689194,-0.00741563543535884,-0.0187007237741963,0.00186122336497685,0.00292643261337266,-0.0141100347452309,-0.00161014140994853,0.00810992836016666,0.0115979115668692
"3005",0.00189688844276836,-0.00774218998111909,-0.00765784318864182,-0.010531709227814,0.00413819916440228,0.000583464961622315,-0.00562689985075671,-0.00833338905612746,-0.00347189443549467,-0.0159236109303792
"3006",0.000227173293111171,0.00352371221984749,-0.000752832345759069,0.00760266234810514,-0.000168067448010678,-0.00252707993104107,0.000738075551883766,0.00135529790083266,-0.00118965839564922,0.00582522978331501
"3007",0.00503537490373973,0.0175569834965958,0.012054954591435,0.0163481719289642,-0.00445821964812343,-0.00272860621743398,-0.016471968300696,0.00730932804254802,0.00212693549321985,-0.00321752554992527
"3008",-0.000339089569466045,-0.00172537721606758,-0.00297783612273284,-0.000247438493297225,-0.00236598289140799,0.000586361986347095,0.00599927364427888,-0.00322494057632128,-0.00220733506912862,0.0129115793058858
"3009",-0.0184646188030989,-0.0143210179714212,-0.0113870298278249,-0.0141089586810673,0.00347259663964605,0.00156243175689497,-0.00198783663122415,-0.00350505697756731,-0.00399898752658046,-0.0152963551974954
"3010",-0.0196184817149225,-0.00926839021465431,-0.00793042491497664,-0.00928956466038244,0.00582362762750366,0.00292514075833727,-0.0369155609639006,-0.00730515978921042,0.00691957127831144,-0.01165045956663
"3011",-0.00109646270673258,0.000407436689290774,0.00278115888932651,0.00679093340357384,0.00598876360343659,0.00246470973809254,0.00897148921382129,0.00109018516962167,0.00237548988609082,-0.0209561733922374
"3012",-0.0149757751750131,-0.00687370337479176,-0.0147283796344791,-0.0166070966735639,0.0132108863931537,0.00349860565428273,-0.0109536414755494,-0.00490070436185508,-0.00609396519519312,0.00401346090748089
"3013",-0.0162779167708219,-0.00410153153879744,-0.00524157361395283,0.00779414682300961,-0.00363112431535351,-0.0012589652738848,-0.0145928083838621,0.00136799735965232,0.0154134207613046,-0.0093271930529496
"3014",-0.0204895814778688,-0.0123552435510439,-0.0308353699995293,-0.00696042806627306,-0.000165565255215383,0.000872740434151753,-0.0124289034106163,-0.0191254622363006,-0.00436092761423901,-0.00874238444107645
"3015",-0.0264228699806871,-0.0125097244568914,-0.0108739256107269,-0.00934587853935331,0.00497017005789036,0.00251883674338327,-0.0360155267403074,-0.00725833723602587,0.0109501009859325,-0.0110645613123692
"3016",0.050524871951892,0.0250725692254563,0.0189332452946753,0.0199161497664258,-0.0107153102153409,-0.00473514613592718,0.0327777124927762,0.0187101767774047,-0.00299944183468026,0.0222376880571071
"3017",0.00767736146002385,-0.00411945709985773,0.0133866627396142,-0.00128469012377297,0.000166558443599918,0.00252431271720477,0.0016137759668855,-0.00367339971543457,0.00760484681247364,-0.00951735773123952
"3018",-0.00129009746574282,0.0085315438866238,0.00118288726889437,0.00951889343605172,0.00841387199929855,0.00542380986725366,0.0030881714297688,0.00226896921766118,0.00406401260678435,-0.00823610138714159
"3019",0.00875894169726044,0.00281966718990634,-0.0017723149860307,-0.00458710591541012,0.00379997008628208,0.00375682634663033,0.00307855345898744,0,0.00156948623111663,0.00276814258750346
"3020",0.0010402261394924,-0.00536804788764733,0.00690470967218171,0.00256017091975935,0.0052671506548716,0.00211130810928095,-0.0216172022825952,0,0.000659810309278308,0.00276057124542151
"3021",-0.0238626985294362,-0.00719598153707024,-0.00568181045197358,-0.0181307745701782,0.0113794138680705,0.00794883503344801,0.00641013602530238,0,0.00906616650348369,0.00825877456338286
"3022",0.0334957623749805,0.0300284400703017,0.0338915979776644,0.0322495719599736,-0.0115751964078068,-0.00807607165956248,0.0107060829555177,0.0209394166858898,-0.00808623703340683,0.0136518996195234
"3023",0.00788462670803924,0.00150783918234376,0.00247757272876825,0.00226770469680582,-0.0029481174909709,-0.00277791840409358,0.0100563706932848,0.00277155517889516,0.00345848973223828,0.00740742970686781
"3024",0.00939531445119868,0.00727724970521004,0.0047528428163377,0.00377064596048715,-0.00262831615057224,-0.00249723574839955,0.0181865305492142,0.00801570574306365,-0.00270804199320496,0.0100266691442319
"3025",0.00467346197184537,0.0122074003189594,0.00548729816065374,0.0177811469305245,-0.00156479460636549,0.000577842414765106,-0.00130374694352309,0.00740325839322598,0.00641816017788321,0.0198544006138881
"3026",0.00352763825236568,0.00147669096411773,0.00602180365869343,0.00713586712479963,-0.00643352333995706,-0.000481357432887575,0.013838205912865,0.00653234675191761,-0.0058866978315214,-0.00259576096476599
"3027",0.000386229700673146,-0.00466944530759072,-0.0115974239925136,-0.0048864049641304,0.00390176191093761,0.0029848359670106,0.00347654100398742,0.00216343551788145,0.00172717334409644,-0.00325304643822777
"3028",-0.00610082392828548,-0.0041974389264956,-0.00359572985025491,-0.00834769879111852,-0.00372096110546538,-0.000576067361145238,-0.00320783086471099,-0.000269926691871536,0.00238089485104531,-0.00848568371229008
"3029",0.011460620413275,0.00223148755734504,0.0121556742124851,0.00693236750180493,-0.00365222095276319,-0.000960423088513185,0.00991224647392364,0,-0.00172003445720481,0.00790000123072776
"3030",0.00241979565566441,0.000247393852239819,0.00487893649240645,0.0122941095971385,0.000999586239192274,-0.000576874772625691,0.00624614084784203,0.00296899300035181,0.00319986880209711,0.00522536480298497
"3031",0.0075868013308118,0.00519411371772183,-0.00205417860801149,0.00437216802979878,0.000249674786201304,-0.00182766858411609,0.00532050651817273,0.00376739364272849,-0.00130854669113967,0.00064975053065397
"3032",0.0133100517690041,0.0125493199315001,0.0132859960627645,0.00483677285386119,-0.00524150296363124,-0.00318051958005638,0.00378024710138813,0.00294900593300329,-0.00892641054027998,0.0103896539161537
"3033",-0.0135105251302371,-0.0133657815503351,-0.0179132240522069,-0.0173285282966976,0.00677479034312034,0.00348060855634302,-0.00288726792138505,-0.00534598377239481,0.0035531318018458,-0.00706942989049986
"3034",0.00209243138848869,0.00689662227975751,-0.00282057702270355,0.010286643122537,-0.000415586253578404,-0.000481687119494256,0,0.00618099784110204,-0.00139973655166081,-0.00129445445557619
"3035",0.000531458931823492,0,0.00584572178549769,0.00969699582542582,0.00656585595161929,0.00318097501064885,0.00352509698584491,0.000801357085242316,-0.00156664744035828,0.00259226447945782
"3036",0.00846143228688123,0.0102738747925124,0.0108736453817031,0.0132052185149609,-0.0047891057586904,-0.00230610966664291,0.0116672426789197,0.0122765386007797,0.014617268630515,0.00517138674472584
"3037",-0.00760012356811146,-0.0046004528226361,-0.00723295343790142,-0.0104266858228054,-0.000995454560206999,0.000288824004975874,0.00905260680336495,0.00580004790948285,0.00349991857805709,-0.0135048870193266
"3038",-0.00132711970563282,0.003162290736064,0.000934134022908761,0.00167640775962075,0.00506590698014953,0.0028887073970445,0.00798819632024106,0.0104849743681636,0.00559657713037076,0.00977835680421557
"3039",0.015830811172781,0.0106692401026993,0.0111981176267182,0.021754736295968,-0.000743582858551251,0.00230404796567218,0.00792487815249099,0.00804167154096946,0.00572672191337187,0.00710137726681648
"3040",0.00878233392598005,-0.00143966380757565,0.00184572243727787,0.00842295418453354,0.00859997491641451,0.00459748344908895,0.010523824154167,-0.00205877078090211,0.000481177312035008,-0.00512816137458549
"3041",0.000481757061891797,0.00120137918419716,-0.00405301062406771,-0.00788867204345278,-0.00603960795429259,-0.00535053761542947,-0.00682312765520365,-0.00128935108379424,-0.00200400801603207,0.00902057392904099
"3042",0.00703533939619638,0.0028799444735339,0.00221968500880565,0.00163710633152436,-0.00446426560040336,-0.00220954597079059,0.00674936576108198,0.00206568145082642,-0.00433735742971886,0.000638547936024469
"3043",0.0041919870151681,0.00909294683762041,0.00406056674540456,0.0137753520561579,0.0045672957539058,0.00173315844328847,0.00610574319325896,0.00154588448043236,0.00258147791692065,-0.00446711284627554
"3044",-0.00131828497181685,-0.00450556635467447,-0.00827202052250664,-0.0135881702274754,0.000495929244277438,0.000768734059336751,-0.00690154771395413,-0.00617438702480122,-0.00675890736046758,0.00128200777892928
"3045",-0.00953282957365598,-0.0131014247312681,-0.013901771695415,-0.0100396617338997,0.00660993328989723,0.00326527490782147,0.00766831447088134,-0.00310640173784338,0.00243029808116813,-0.00960307277514072
"3046",0.00122153479240406,-0.0036205910115541,-0.00883458626411948,-0.00566050925359562,0.0042682938621712,0.00133997641522599,0.000237945840694032,-0.00103865603094089,0.00379829487309347,0.00129284668618146
"3047",0.000554490663109197,-0.00242247318635835,0.000948170757803402,-0.00332061446599796,-0.00392315371120699,-0.00152947231739975,0.00285296522423062,-0.00285951521082994,-0.00491104584905433,-0.00581019987504727
"3048",0.0128595385404742,0.0109276137047758,0.0176203108923771,0.00832939014270906,-0.00254361825249771,-0.00134037007979548,-0.00580845712218381,-0.000521358812938466,0.00210358417643342,0.00584415558710938
"3049",0.00324681406465155,0,0.00242046825771447,-0.00708050100986224,-0.00378424305713032,-0.00249244999892939,0.00465010208765881,-0.00756388830315857,-0.00395606326533127,0.00581019987504727
"3050",-0.00221803740926252,0.00024020320625362,-0.000742962608969666,0.00190163700867041,0.00569779580830776,0.00470913807536011,0.00320432526948089,-0.00289096435785263,0.00559289116658279,0.0025673722456947
"3051",0.0108972347563729,0.0158500759443467,0.0128252875808565,-0.00142356956944245,0.0015601086842576,-0.000956323283694771,0.00615172616715309,0.00711638876670939,0.00596489611421736,0.0185659623806202
"3052",0.00173039075714576,0.00401902024241663,0.00165172024661309,0.00784030552574144,0.00254119836673117,0.00172332708772571,0.000235093807417375,0.00366398180854843,0.0152243105314669,0.00251418451559937
"3053",0.00201546881511128,0.00565095250040581,0.0010992312621565,0.00565774417866449,-0.00286198379442271,-0.000191270735674043,-0.00705292803421931,-0.00260753099905153,-0.00173633784695348,0.00313475350515446
"3054",-0.0035557463812157,-0.00468270588283959,-0.00146411335623353,-0.00210963338775172,-0.0089386851112796,-0.00296360788603089,0.000828630872581115,-0.000522829622447096,-0.0113061350891966,0.00312495753357278
"3055",0.00620003789330359,0.00305814574866936,0.00219941826476155,0.0110406305881516,0.0059576617418442,0.00297241696438721,0.00532278492743155,0.0031388186823178,0.00359853649903541,0.00249225404025921
"3056",0.00136116290080412,0.00211069496809646,0.00566939857034465,0.0111523657784109,-0.00296128601272005,-0.0015293841314572,-0.00729482750364208,0.00104307505532364,-0.00103583266932272,-0.014916033180699
"3057",-0.00071542406777203,0.00725489906385612,0.00345516241274413,-0.0034466771954148,0.00495014108910796,0.00296792231409171,-0.00272607246368051,0.00442841421688955,0.00167503385957479,0.0044163819462697
"3058",-0.000429604075305234,-0.00348525128702581,-0.00525561257196572,-0.00853122863455436,-0.0113291111173774,-0.00353216194086881,-0.00285239766452616,-0.00440888982650112,-0.00708711566989773,0.00502508265366841
"3059",-0.00186260875154964,0.000932658895962613,-0.00965560334517146,-0.0130232728235646,-0.0034043388399102,-0.00258681484711731,0.00297975826807462,-0.00468879034944547,-0.00561395451737989,-0.00250004222829769
"3060",0.00624397335399918,0.00628940702111547,0.00294329064045051,0.00117813712716908,-0.00924304773938445,-0.00328139886960854,-0.00213903786607894,0.00209379372670249,-0.0170175097510687,-0.0112781954887218
"3061",-0.00363759523044205,-0.00416666796219789,-0.00311812862311955,0.00141208152733818,0.00783747766496079,0.00308960364550814,0.0041681445294075,-0.00365629769116516,-0.002625525171288,0.00316865365604024
"3062",-0.00136000950695603,0.002091954792103,0.000919984011975794,0.00987080186106781,0.00209055898253485,0.000577554423839333,0.00308342547166962,0.00550458720849401,0.00131624714241929,0.00505365229360066
"3063",-0.00605693835380283,-0.00185572667612555,-0.00588232820768719,-0.00558539840574235,0.00367147177326399,0.00278984613651945,-0.00484736980387412,-0.00599592530939208,-0.000903713433259012,-0.00565681936947671
"3064",-0.00836548785064783,-0.014640834209391,-0.0118344016466634,-0.0184880609159473,0.00648481942829515,0.00335755297243434,-0.00178234298268354,-0.00131098712506839,-0.000822292567862037,-0.00252848771387459
"3065",-0.00199998717299044,0.000707523013688149,-0.00168415460981863,-0.00715319349546928,0.00421293196230077,0.00143414444343404,0.000952272023947209,0.00709002324085284,0.0109455516262769,-0.000633692099297978
"3066",0.0145013186024046,0.00848454121261688,0.010871684599586,0.0187319824896492,-0.00296133309895363,-0.00076362198711788,0.0147443329811174,0.00547610844061741,-0.00488438635247102,0.00126825226655392
"3067",0.00377101020321624,-0.000934838417954387,0.00241057528928112,0.00518630593197988,0.00701255423388281,0.00277076398027476,0.00410132867402768,0.00233398818279862,0.00605370592365362,0.00633316485474422
"3068",0.00661917441811677,0.0109941885240021,0.00388454321044551,0.00117261114028877,-0.00188429746418195,-0.000380969249435537,0.00455124033133969,0.00569208527816278,0.00699294990259514,0.00629318041424543
"3069",-0.00063972682814073,0.00439610648327671,-0.0106873085292396,-0.00538763571787149,-0.00722319600732779,-0.00142999325654802,0.00151023877279588,0,-0.011547093396224,-0.00437765136383261
"3070",0.0049404793267831,0.0110573163994638,0.0115477232206478,0.0146020521884305,0.00661441822819397,0.00315001335426235,-0.00231985586903449,0.00514529442180911,0.0045747649840775,0
"3071",0.00362581486188995,0.00455690341593651,0.0027619472276974,0.0111419380421767,-0.000574929191366924,-0.0013321158919477,-0.00558083549199873,0.00295669084999695,0.000569244526557489,0.00502508265366841
"3072",0.000248042021727013,0.00362895767333882,0.000367224067863603,0.00045919480299994,-0.00221885971106273,-0.000667131016361733,-0.00292288679397656,0.00179455020211283,0.0027632964664881,0.00250010572949733
"3073",-0.0030099613115413,0.000225887591245533,0.000550624524082055,0.00160630244880355,0.0104603543386219,0.00696040526398689,0.00334210767114684,0.00614110584811067,0.00648405754135339,0.00748116896669782
"3074",0.0112947065122899,-0.00271113613143625,0.00660436383577889,0.00137446093798088,0.00220089812115432,-0.000473334533592107,0.0169491488620348,-0.000762887181214089,-0.00402641327105813,-0.00495051590324702
"3075",-0.0192464328787829,-0.022881754862752,-0.0107526929746663,-0.0292839178927583,0.0155346253251736,0.00738918292998458,-0.00601847966956648,-0.0106898200425055,0.00234476875808531,-0.00870642553817436
"3076",-0.000751999205660159,-0.000463794358181224,0.000552653338020903,0.00235682954229377,0.00160181354547784,0.00253897185525975,0.000232822368848806,0.00643174828237369,0.00766312004788983,0.00376411527292286
"3077",0.00745419071814113,0.00417543894801375,0.0110477513066725,0.00305661626897291,-0.000719491264476346,-0.000844228428811933,0.00745051448102241,0.00408997739022321,-0.00496313648676172,0.0018750634218232
"3078",-0.00522907918056825,0.00207900277369832,-0.0034601964802311,-0.0107828494197302,0.00920215752647913,0.00291039960286965,-0.0020798945453756,0.00127296711619262,-0.00522929190918853,-0.00561453565263736
"3079",0.00379048034988494,-0.00437996354663039,0.000548209468230754,0.006635030683249,0.00348859816728653,0.0000935877008350072,0.00868452505655792,0,-0.014152850559598,-0.00313672023395206
"3080",0.00630541454698763,0.00463066352589037,-0.000547909099274824,0.0103577666242571,-0.000948150988453023,-0.00159131927973732,-0.000803578085584622,-0.0012713487310646,0.000902378984374508,0.00062924131247688
"3081",0.0118591013133493,0.0124453407572034,0.012609657522384,0.0165424079595653,-0.0142037948935785,-0.00687634768193757,-0.000344702900577087,0.00305496052894005,-0.00393412828564654,0.00943396226415083
"3082",0.000489899471532551,0.00318692074067584,-0.00685805625158564,-0.00320873483896256,0.00184916948980818,0.0017027147133073,0.0064360485909154,-0.00456852564940724,0.00370282237885977,0.00249225404025921
"3083",0.00157355791258795,0.00816880156406663,0.00599674240995562,0.00689815647109082,-0.00866775529817598,-0.0031161836471818,-0.00102767443561325,0.00382457738773323,-0.00147565170989539,0.00124302907589291
"3084",0.00265349720121977,-0.00135055564056674,-0.000541871823048989,0.00616577051179457,0.00283363990284746,0.0010418784668309,-0.00148610581393005,-0.00482603487065947,0.00254513951038238,0.000620774470232011
"3085",0.00484028262048652,0.00157765881058602,0.000722899780049913,0.00771678980591073,0.00129160104824799,0.000473219539410152,0.00686895783834607,-0.0076569364766691,-0.00106459748534438,0.00310163159940502
"3086",0.000762254906854887,0.00180028157779355,-0.00234777321903079,0,-0.00354742190107149,-0.00160781001581611,-0.00591249351119671,0.00282927261442301,0.00434496628107151,0.00371063797274185
"3087",-0.00512482914563506,-0.00539086066455974,-0.00543089582866263,-0.00202705106742251,0.003155557061292,0.00179973830349667,-0.00480386850924797,-0.00641184113733062,0.00522406325648417,-0.00184842871977575
"3088",0.00341109415008267,0.00338755847421179,0.000181998558285823,0.00473933087900114,0.0024197154007346,0.00236420436039064,0.00907941117720523,0.00877645302167895,0.00308564347404561,0.00864193295515259
"3089",-0.000277599964199959,0.000224972454013761,-0.00309372840647026,-0.0107817377047476,-0.00587389290150764,-0.00226421229530682,-0.0010249823619034,-0.0033265911555368,-0.012790431577677,-0.00489591927758426
"3090",0.00676597042441673,0.00630078789608879,0.00511136584719796,0.00726619820166841,-0.00712241614409814,-0.0046332638632276,0.00524453226761756,-0.000513478546651958,-0.000983968863894291,0.00307492641515528
"3091",-0.000654799203336998,0.000894331420260075,-0.000181601905736906,-0.0051849025071149,0.00252695111999879,0.00133013675655835,-0.00510383526358982,-0.00410993873858567,-0.00188790935093308,-0.0018393001365179
"3092",0.000655228246270623,0.000223498496151997,0.00399637568647071,0.00747787103855768,-0.00626110372603317,-0.00341528957280846,-0.0214317803771086,0.000773709622975627,-0.00896378304216749,-0.00368550360883424
"3093",-0.00244697931209048,0.00402052772631456,0,0.00292402188840568,0.000409128171228401,0.000190316421467607,-0.0090866441350117,-0.00541231266030817,-0.00190858016913809,-0.00369913679082623
"3094",0.001969209231794,-0.0020022253998031,0.00144742452087487,-0.000672835386063775,0.0052346805745338,0.00237959226801587,0.00681873366918651,0.00155486250818893,0.00074828733578558,0.00309401742611271
"3095",0.000861989469204349,0.000445816278181077,-0.00361334050228201,-0.00650811577890575,-0.00480072295598799,-0.00142447224296738,-0.00980854010239374,-0.00155244866396542,0,0.00493537152270385
"3096",0.00899165105234245,-0.000445617614594718,0.00562100869055659,0.0022588724872199,0.00212585414467625,0.00180678991874017,0.0119104327278994,0,-0.00207692941571169,0.00122758060901673
"3097",-0.00221929290105549,-0.00557288773693843,-0.0122611159378654,-0.0135225033359181,0.00815856399607062,0.00379636508195302,0.00652604018357827,0.00207304669904329,0.00291373619096569,-0.00367860027303579
"3098",-0.00061615100889556,-0.00201748556978421,0.00219064128530899,-0.00137088085325665,-0.0014567058238163,-0.00122913213284936,-0.00196827896603968,-0.000775710466209167,0.000830073870423442,-0.00184621621650349
"3099",0.00465695313555914,0.00134763973897556,0.00910750637412527,0.00388933748492981,0.00340386439451823,0.00265070544861867,0.0075405215300397,0.00258804654094003,0.00663517458737672,-0.01171384965108
"3100",0.00156763398292603,0.00471068089012761,0.00397107225475857,0.0020509788130334,-0.00638073610962808,-0.0020772117073482,-0.00955665264832328,-0.00154881389422157,-0.00444921303989754,0.00062387250715612
"3101",0.000510523581929156,0.00468852521263408,-0.00359587334694511,-0.000909732416538689,0.00512118599939471,0.00198698721349788,0.0113927195504564,-0.0025853982135331,0.00306211200757911,0.00311710095042761
"3102",-0.00751643657449186,-0.00755557381194549,-0.00342835436595113,-0.00751191561836884,0.00412500493812895,-0.000454352153353765,-0.000689722735418674,-0.00285118861810774,-0.00660061897526276,-0.0031074148247241
"3103",-0.00215899961987986,-0.00425433721474,0.000362104342996439,0.00229358431583759,-0.0047618436953536,-0.0028396770015352,0.000345099390604897,-0.0122172773666047,-0.00382059794317935,-0.0112220701642258
"3104",0.00978776365603973,0.00966952893446882,0.0128507441983778,0.0118994028090658,0.00283843842797782,0.00132902132890256,0.00793373464372582,0.0202631176853336,0.0059196263811967,0.000630495656581909
"3105",-0.00411524659860074,-0.00913143646228798,-0.0101858689660194,-0.0205789598319196,0.00274940151337888,0.0025597560465509,-0.00330819824749007,-0.00412690004495075,0.00132611684498762,0.00315068397557128
"3106",-0.016699636164017,-0.0188806534752602,-0.0182343226885366,-0.0196259817452258,0.00766124746571606,0.00340423627385533,-0.0181984549139697,-0.00207194464060401,0.00331099252232425,-0.0125628342747678
"3107",-0.00138930551079675,0.00504003807611109,-0.00606843938505597,-0.0014130791503687,-0.00432170332776405,-0.00188497487607886,-0.00011658871364606,-0.00285511409253092,-0.00247500208295515,0.00127222146063866
"3108",-0.00302581413683745,-0.00569867301107108,-0.00647540539013314,-0.0158018909141748,0.00409939203447029,0.00264389106393192,0.00233186692208909,-0.000260167797899835,0.00239842023328363,-0.00508254897919436
"3109",0.00502348253674034,0.0066483844030798,0.00689003080324002,0.00599081150444158,-0.00136086348109921,-0.000659229834115482,0.0105850278208577,0.00702950076424536,0.00189771456842536,0.00191564380807363
"3110",-0.0251302685601803,-0.0214074238214267,-0.0225633558986281,-0.0333491113189348,0.00785566532681647,0.00499436355348482,-0.00115104312184344,-0.00646334092660938,0.010211628098493,-0.00509874586703907
"3111",0.00904367806562911,0.00791249180288123,0.0140020005452519,0.014046325565674,-0.00294286077225636,-0.000937572517234364,0.00414847368639659,0.00468383823151197,-0.00171190187840398,0.0134529142144599
"3112",0.00585742906501041,0.00600314713556593,0.00149270465324158,0.00194405215377813,0.00614244982433032,0.00319083342969662,0.00654120389075019,0.000518000240836036,-0.000571615225964495,0.00884951432741188
"3113",0.00926133772193305,0.00895116447166222,0.0040992095080199,-0.00485085013684705,-0.00332996564858268,-0.00196451968126155,0.00592857832361804,0.00569499631699255,-0.00719010545951559,0.00563909774436078
"3114",-0.00646503774102314,-0.00636942136213858,-0.00371129058040376,-0.0180355533973179,0.00222729168406333,0.000468654412589142,-0.0028335139367841,-0.00669237552085244,-0.00707760666484059,-0.00934579439252337
"3115",-0.00661216256784525,-0.00663925184619996,-0.00540138999392958,-0.0042194821409961,-0.00206362279503691,-0.00168642265985042,-0.0147760080709701,0.00492358100411305,-0.0000829092402335752,0.00440255832365777
"3116",0.00901569426577886,0.00691408613603706,0.00692881581097637,0.012711982230929,-0.0015906349038487,-0.00112622865174539,0.00842169582992347,0.00360999422839448,-0.00232093834815106,0.000626152843005601
"3117",-0.00307148747575614,-0.00389105996974504,-0.0081829627278277,-0.00492258566601023,0.00573560320029465,0.00300658625004013,0.00354648921639433,-0.0069371647045674,-0.000997033890021259,-0.0143929485468923
"3118",-0.01221855881842,-0.0101101873239111,-0.00750040841760746,-0.0128617317508564,0.0112473870545446,0.00608900728374207,0.0013680414172963,-0.000776224331982656,0.00773453106677535,-0.0209523796007606
"3119",0.00226843873144689,0.0106776838857965,0.0154920762800805,0.00100238166212985,0.000861786816457988,-0.00027929810817473,0.00330141906729553,0.00828585781520452,0.00107291410535471,0.0136186761454711
"3120",-0.00930064308716261,-0.010564875485074,-0.0083721113143046,0.00350430742940389,0.00719984403007801,0.00437725858565852,-0.0105525575108755,-0.0118130115214424,-0.00387469899732817,0.00831731624288978
"3121",-0.00671065758038458,-0.009285165666017,-0.00469040353701378,0.00648540514297902,0.00303031760173256,-0.000370843553664013,-0.0119265991102806,-0.00077965359554466,0.000331051885607003,-0.00380710643535986
"3122",0.00273121289952494,0.00585753881111506,0.00452402452182943,0.00545226665115939,0.00859859142780106,0.00361768549343844,0.00406223920630433,-0.00182048862857032,0.00678413981672543,-0.0101910607913405
"3123",-0.0134754076712191,-0.00931751345180587,-0.0106961373725604,0.0034508556212296,0.0125191323056515,0.00665514810979939,0.00416132615001774,0.000260467225622119,0.013476867228583,-0.0263835464521808
"3124",-0.00254290553998304,0.00705399313841748,0.00588009518602739,0.00908876167101114,0.00668912388103027,0.00481149173029927,0.00391391221824744,0.00859598415636453,0.0144328141663372,-0.0033047148998443
"3125",0.0217067691661179,0.0121408250304145,0.0115028899140681,0.00219067259089889,-0.0114014127826573,-0.00366244594942011,-0.00321068532849922,0.004132229316262,0.000319726638000839,0.00596816962723756
"3126",0.00866210017382674,0,0.000559247266923357,-0.00801550806780282,-0.0056519719533592,0,0.0209363632790209,-0.00411522426590738,0.00255692365070836,-0.0204350464341544
"3127",0.00650265505545078,0.00553645399280267,0.00111802157860419,0.000489777815857018,0.00322611386254312,-0.00018357420286419,0.00146483999458713,0.00335740823809583,0.00326768149145074,0.0174966572558402
"3128",0.0100070266830656,0.0126176168298731,0.0120975126305463,0.0078316013284323,0.0086515869319348,0.00395216791774766,0.00303774406368307,0.00566283095592479,0.00564028453225962,0.00330683328664261
"3129",0.0045890253470533,0.00203887392717506,0.00459726956093376,0.0104420309138338,-0.0094123577801335,-0.00494370754001927,-0.00302854412175546,0.000256062048445971,-0.00995334576043438,-0.00263676074053543
"3130",-0.000242233605321607,0.00520012368932532,0.00329488136825185,0.0112953525142874,0.000613096679436875,0,0.00168766121601283,0.00511762066655463,-0.00119685628027033,0.00660936264706513
"3131",-0.00176527846676466,-0.00584796313740699,-0.0111293988469486,-0.0106939452238819,0.000765718471174015,0.00257599416888787,0.00325729141732722,-0.00865579992822318,0.00519253874420822,-0.0137885081622434
"3132",0.00412615805111671,0.000905040058121198,-0.00110693817028551,-0.00168144473718868,0.00344364856424706,0.00247782169812183,0.00369458786589671,0.00308163454097854,0.0061193355142759,0.0126497765772546
"3133",-0.00110491755873576,-0.00791147278110738,-0.00258585627527896,-0.0110684439992836,0.00251660395058506,0.00073224373888725,0.0016731660306013,-0.00409614876056053,-0.000315955771184151,0.00394477291203388
"3134",0.000380167479839155,-0.000467698857587906,0.00293375329657919,0.00394719683044364,0.00174957024357814,-0.000182799489711782,0.0107165461696976,0.000513942841349424,-0.000632071754615549,-0.00458419598484128
"3135",0.01047111872822,0.0142722553725101,0.00596243420023201,0.0241758211060821,0.00501156548636028,0.00192119235623034,-0.00177637704113398,0.00668042306440619,0.00506008843152861,0.0118421049993025
"3136",0.00225713436313479,0.00438300432490513,0.00889057583554731,0.00834530156760138,0.00143566485670354,0.00273954903834883,0.00622849106778434,0.00280763680541285,0.00605723711318662,-0.00195051907153276
"3137",0.00955436453849523,0.0101056230765517,0.00973010138533414,0.0146606681790564,0.00264080438932068,0.00163922018595719,0.00442134670406569,0.00763549876929681,0.0251779030821637,0.0201954158937032
"3138",-0.00145356932447815,-0.00159161744179992,-0.00981819195421363,-0.00326268933584439,-0.0109866616596832,-0.00409131620320091,-0.01265543037629,-0.00303103940568195,0.00663561126812895,0.00255425662399422
"3139",-0.00122451041173965,0.00159415472626723,0,-0.00140287256701155,0.00745651416551274,0.00346917571314931,-0.00624160151638264,-0.000281951425623261,0.0148507808713678,0.00445857696222429
"3140",-0.00980788024558843,-0.00568439378333985,-0.00440685919472805,-0.0103020413273999,0.00309652912349612,0.00154653121802184,-0.012786139150528,0.00102520383934634,0.00194113032789112,0.00317059845271306
"3141",-0.000997519241488276,0,-0.00147551117842637,0.00946294278569781,-0.00639986445630936,-0.00408772861193096,-0.018859244880739,-0.00512030139991004,-0.00916539513782555,0.0050568469803165
"3142",0.00354602859561637,0.000228765869366043,0.00406355357645305,0.00703082580433767,0.00704723862168843,0.0030099124245051,0.0115793832379076,-0.00257349292328179,-0.000977701729880986,0
"3143",0.0051457252016176,0.00754453222843843,0.00404710793652341,-0.0013963429297108,-0.000677371672561877,0.000454657006253134,-0.000572388366601229,-0.000257902326172399,0.00271003470972686,-0.0106917812989837
"3144",0.00907863161519162,0.00294984718437985,0.0142909140502754,0.0118852969304599,-0.00233864786733473,-0.00125637233900422,0.00343601751777167,0.00335487152695868,-0.0193693848206319,-0.000635706350688436
"3145",0.00260428934286128,0.00316739058927706,0.00307079620621087,-0.00253331342675633,0.00771310523278301,0.00355551717066671,0.0156375091020537,0.00488681722784201,0.0213597389894249,-0.0165393960464058
"3146",0.00799514606070084,0.00721693661030542,0.00288129605840015,-0.00184724552277449,0.00712891326403531,0.00190761456814914,0.013261474736179,0.0133094644502609,0.00164905924146463,0.00970239117406657
"3147",-0.00113792097386289,-0.0107478835265966,-0.00430952706425625,-0.00693958302491282,-0.0132625874675875,-0.00634692946889814,-0.00454756375903886,0.00176806528259421,-0.0111502353083054,0.00192190997549258
"3148",-0.00549479412677034,-0.00452691514113779,-0.00577096070937277,-0.00605645743371463,0.00135909457122119,-0.0010037182904411,0.00323133103173867,-0.00353002504447941,-0.00643261697012709,-0.00127885885720846
"3149",0.00124650819394789,-0.00409277634153993,-0.00888806542699261,-0.0030465611281224,-0.000377017270022373,-0.000639458116921343,0.0048867176921128,-0.00328939716477317,0.00350374761616434,0.00320104594039505
"3150",0.00477797848780703,0.00365300231091514,0.00603956233632985,0.00846262446303525,-0.00550689835262541,0.000548554124587985,0.0053048811023475,0.00203092912728287,0.0157874914611007,0.0216975534556096
"3151",0.00234424810568612,-0.00159241021582646,0.00181915544171485,-0.00186482854745662,-0.0133505335560106,-0.00493293082051971,-0.011213638246575,-0.000253344791419141,-0.00844358501914999,0.000624588412292182
"3152",0.0044769180542914,-0.000455657414430433,0.000363170424888093,0.000700641088742904,0.00115327135730303,0.00110158956018158,-0.00177894459939676,0.000760335966915715,0.00625472508488456,0.00249679418045523
"3153",0.000332638466449042,0.00182362115195867,0.000726058791346462,0.00373386604585724,0.00575933279631768,0.00210920514445179,0,-0.0020258678313535,0,-0.0105851998891362
"3154",-0.00322526608279028,-0.00341302830231749,-0.00743696469138722,-0.00139494950010655,-0.00297738981738749,-0.00219625235539789,-0.00233906331001332,-0.00304495681329786,-0.00846255529440998,-0.0106985729502709
"3155",-0.00680500124659,-0.00205482098192666,-0.000913770348274223,-0.0030267948703101,0.0107978018738566,0.00467724616463361,-0.00401917374946337,0,0.0164653179667065,-0.00890587338578497
"3156",0.00366091494574561,0.00503319463611973,-0.00256079339209137,0.00607203990052496,0.0000757100139177069,0.00246455808173129,0.000224154913402552,0.00432681148081171,0.014117951937614,-0.00706035519196246
"3157",-0.00555490281760429,-0.00614610619737521,0.00256736789082113,-0.00510682702313581,-0.00234863761284743,-0.00182109430722421,-0.014681210267398,-0.00405476184650233,-0.0147273963870866,0.00581777724944499
"3158",0.00245638302451745,0.00206134073216435,0.00146338454895445,0.000233249618771136,0.00189862533345653,0.000456014182742548,-0.00181980514145208,-0.00559783192458008,-0.000148761804500963,-0.00321338909511093
"3159",0.00715004130034846,0.00640005437435875,0.00803648435627458,0.00116630967482623,-0.00545715146052583,-0.00164126263003339,0.0101413078418933,0.000511553451062463,-0.0056526219186156,0.0064474309978213
"3160",0.00469958129466197,-0.000681415714134492,0.00126829611388213,0.00163101228300588,0.004343699410021,0.00146133853893038,0.00282011243001823,0.00153470066860928,0.00508634146029863,-0.00448428304224902
"3161",-0.0047770471638533,-0.0104544921902794,-0.010676765512232,-0.00883931988352438,-0.00478022440332493,-0.00173267521354181,-0.00461201744467032,-0.00561806375548102,-0.00707000844943095,-0.00386106898946703
"3162",0.00669998378280923,0.00528251789330536,0.00256084892148234,0.00211223448544939,0.00236367169984364,-0.00018288491538454,0.00339029080426023,0.000513613590390705,0.00164893571651836,0.00129201154218861
"3163",-0.00182115423070373,0.00182771844773733,-0.00127714463139084,-0.00187356305370401,0.000304045582917079,0.000913815157803421,0.00292831346862665,-0.00359333909634241,0.00665968277955487,0.00387103320698201
"3164",-0.00245474523732159,-0.0150513285907889,-0.0063938890780636,-0.00774281072390437,0.00243337525264486,0.000456421147537744,0.00718687290381648,-0.00644005679095649,0.00334495654013933,0.00578399589622292
"3165",-0.010940395706309,-0.00648294383027359,-0.000735421822407156,-0.0122960575234992,0.00804066243010082,0.00255503428485171,-0.00334483985762701,-0.0111484985459063,-0.0131129726807816,-0.00638968965774234
"3166",-0.00870786008857782,-0.00419483324743752,-0.000183953528870129,-0.0196313501550002,0.0198602356012916,0.0113424462316467,-0.00100679685157012,-0.000524499541312951,0.0240221967708476,-0.0276527736668752
"3167",-0.00752947380429148,-0.0100632799074319,-0.00515274518193776,-0.0097680498451983,0.00924154683514855,0.00207367280733006,0.00447926352014805,0.00996852084646327,-0.0038120737830929,0.00132277363287803
"3168",-0.030073177128459,-0.0217492986935625,-0.0247872446882911,-0.0369913456359242,0.0172880869670258,0.00863688972330068,-0.0179487523718886,-0.0199999603426408,0.0139818530722045,-0.00858656973011873
"3169",0.0140229710656532,0.00410817693262899,0.0127085959851618,0.0143406376016595,0.00799308291406065,0.00160552677761361,0.0105574192384557,0.00477073795400651,0.00812839144276589,-0.00532973477973142
"3170",0.000590706734606261,0.00505412797474047,0.00693008501657366,0.00454429455290373,0.000357231013315973,0,0.0104470331619766,0.00501185603401866,0.0151896907295461,-0.0127260991363837
"3171",0.0196200432930607,0.0107759048765264,0.00706851242864848,0.0123146483099983,0.00214241113127467,0.0000890839402085675,0.0167872345872235,0.00524943005026923,0.00503468997206946,0.00542736221015194
"3172",-0.00681157174872604,-0.00497507715621748,-0.0105282273865946,-0.0101788182562097,-0.00199535413310803,-0.00151373440370495,-0.000109448131649592,-0.00365548519574965,-0.0033161716874669,0.00877197552943043
"3173",-0.0121732525383303,-0.00785721171229481,-0.00952025085147989,-0.012039095242882,0.0208497890549098,0.00633188534516615,-0.00382716682085837,-0.00445482531172781,0.00969849956457947,-0.00735781389097367
"3174",0.0155516769320576,0.00863932367315479,0.0113078755944878,0.0126936034863279,-0.00342731295926657,-0.0035448790518019,0.00109768998778548,0.00236910024880554,-0.00595951742412126,0.0235847893992234
"3175",-0.0295676050817044,-0.0271235133822006,-0.0242265731886174,-0.028829206667189,0.0225294421678923,0.00667029809802799,-0.016228031964407,-0.0168067597039955,0.00684159265652129,-0.0151414293457932
"3176",0.00264184678190471,-0.000244457787457741,0.00954929276952798,0.00671132039367262,0.0111195849342762,0.00636103568713708,0.0110342458558053,0.00988246217922661,0.00665497022767081,-0.00802138964796029
"3177",0.0147548817774983,0.0119862114749407,0.0104048131904593,0.0138462212519352,-0.00801040970349742,-0.00263374733746802,0.00870910206080366,0.0134884144580947,-0.00640221307729039,-0.000673900029193431
"3178",0.0120477635485325,0.0077350491748287,-0.000187191054237923,0.00404646369744643,-0.0143023839106715,-0.00475312895888846,0.00754100599093888,0.00287059405438028,-0.0116963020849999,0.00472013878150723
"3179",-0.00766242014277529,-0.00575667356436949,-0.0020599419144286,0.00201511649957387,0.0103443749307404,0.00442208547943634,-0.00748456484262106,0.00286237733103234,0.00779537943593356,0.00268454096763349
"3180",0.00813536575527629,0.0118213588260563,0.00337778586630177,0.00955249609479702,-0.00666530946935318,-0.00264157003914878,0.00371576394418005,0.00337304020137297,-0.00316441866147987,0.00334674288307091
"3181",-0.000307831231642131,-0.00214587850316972,-0.00149622642837766,-0.0129482152012312,-0.00664072951795036,-0.00220707179369384,0.00555322264925273,-0.00362028702041883,-0.00253951052975143,-0.00466975715446305
"3182",-0.0256874004775369,-0.0126642052673843,-0.0112380586884105,-0.0148839119335499,0.0164345097063081,0.00672429823982501,-0.0137519807504317,-0.00207626004178918,0.0195898452442651,-0.00737260842225429
"3183",0.0110583387168111,0.00701842345292092,0.0145861004558192,0.00537771948421817,-0.00404219765149383,-0.000966673640810156,0.00735614879041946,0.00520156152270079,0.000138752863130476,-0.000675265120282376
"3184",-0.00392358128106918,0.000480624892194026,-0.00317401585972565,0.00178306281537877,0.0154090161852407,0.00431080359009739,-0.00381474132292792,-0.000517467310621189,0.0095707398630871,0.00675673356420781
"3185",0.00704154482058694,-0.000720699816569192,-0.000374598165568285,0.00279675722004358,0.00128719003474886,0.000350295254418986,0.00229760512883814,0.00232973891320598,-0.00281653486490541,0.00872487747592454
"3186",0.0127730008955875,0.0100961790678529,0.00712008917882345,0.011156294873903,-0.00378881393838737,-0.0019263782405835,0.00796851607087046,0.000516642913496179,-0.00716456993208681,0.00266132126566654
"3187",-0.000444266610053812,0.00356969475049329,0.0031627773106373,0.00777320015145233,0.000271463971838193,0.000263147420931364,0.00129959454927864,0.00438812856130921,-0.00256727041934735,-0.0159256794434508
"3188",-0.00584717438145466,-0.00308265942902075,0.000556411697061998,-0.00622041509891968,0.0012923756493497,0.00219652969625006,0.00973389595621588,-0.00565416056497348,0.0139130434782608,-0.0053944247471307
"3189",0.0113503794815639,0.0164129025794546,0.00556070388652974,0.0167751472495858,0.00149433234096996,0.00157794465322669,0.00781914937773287,0.0129232542012603,0.00624359519725548,0.0237287654582146
"3190",0.0128553428673219,0.00514855841283213,0.00718896000714198,0.0113272456274078,-0.0181101077677718,-0.00805257182616159,-0.00627045670859405,0,-0.0240011243965328,-0.00132452568052432
"3191",0.000772249250603263,0.00209551025870502,0.00347728897432753,0.00438284889779061,0.00711509672066946,0.00061765403531111,0.00192508157137761,-0.000765382299363626,-0.00852313125976756,0.00265256475118081
"3192",0.000503305196656756,0.000464656192306956,0.00656573703473406,0.00315151057762009,-0.0177652006225232,-0.00617287002698497,-0.00651153240588676,-0.00229831752975751,-0.00373449131531134,0.00925928103607609
"3193",-0.000234632340077701,0.00139339129405336,0.00289904636497629,0.000724899529996215,-0.0175279676911486,-0.00727590543585888,-0.0106371625076983,-0.00307142757480161,-0.00855793202176902,0.00131050490558815
"3194",0.0071108336694321,0.00533390108254062,0.00885281146502215,0.00700316587316152,-0.00177685381711112,-0.000983245420517642,0.000977461867549323,-0.000256754661383529,0.00606367557744147,-0.00719890871020412
"3195",0.00346387255822345,0.00599775261627977,0.00662602489682618,0.00719429870050825,-0.00655089160666489,-0.00223660936898373,0.00488230511222287,-0.00154078554687309,0.00205635681809802,-0.00395517459858208
"3196",-0.000663856979901234,0.00275165937693567,0.011741671559945,0.00571429432984538,-0.0213589625401879,-0.00914629641549203,-0.0116606170280036,0.00823047122520904,-0.00827917451207039,0
"3197",-0.00308870394850747,-0.0107477833270933,-0.00527511763671229,-0.00781256309453338,0.0127435919048571,0.00434388645230133,0.0102688007919778,-0.00433685496167135,0.0083482914740618,0.0443414722905136
"3198",0.00253189104649021,0.00485441592267422,0.00371219485965035,0,0.00542359553954452,0.00261296177881887,0.0109212533874659,0.0061492063117754,0.00198131181807826,-0.0190114068441065
"3199",0.000598226077207942,-0.000920212368100692,-0.00211345210204517,-0.00405627178753709,0.00424384090488927,0.000359619249856502,-0.00352976269731375,0.00050927011243207,-0.00628530340599009,-0.00645992644230764
"3200",-0.000066511411233372,0.00345389364657311,0.00741266847814037,-0.00407289001775268,0.00300807673000203,0.000449072551662377,0.00483033402077027,0.00610840432256432,0.00405082774247889,0.00520164843502324
"3201",-0.0047247367713863,-0.00206512466072295,-0.00227751745562499,0.000962295325206863,0.0132106299142039,0.00574718394542972,-0.000427324620401959,-0.000758799181866721,0.0118204842286274,0.0012935513870731
"3202",-0.000234727581092775,-0.00252933908112429,-0.00105352723640928,0.000961345657114476,-0.000211472972139748,0.00142856988504336,0.00149622121804072,0.00104761520820662,0.00559638346826974,0.00258408871869475
"3203",-0.00784682088711497,-0.00576301561431658,0.00140619036464584,-0.0105643026372392,0.0120541737923394,0.00499279451241974,-0.00124672118125113,-0.00357411506328831,0.00528692173913048,-0.0115980023440451
"3204",0.00591481719694231,-0.00486914070573119,0.00403720693090559,-0.000727989074488233,-0.0146271373303023,-0.00656482459099494,0.000753304591408988,0.00358693518235453,-0.0185453815841596,-0.00586701408252943
"3205",-0.00208321803963207,0.0053589206084248,0.00174821624234922,-0.000242864611907589,0.00643260422855896,0.00214316091194666,0.00817200205059088,0.00638249788437895,-0.000282091232008841,0
"3206",-0.0053871747802523,0.000463378343763532,-0.0143105887060947,-0.0128734131819004,0.00245814763670404,0.00142570641567441,-0.00607932131171751,-0.00329778661023139,-0.00514842397939885,-0.0039344926789654
"3207",0.00463772364056836,0.00231654147395277,0.00460340617119259,0.00565945449583971,0.00245221903135873,0.000801007691797029,0.00375572162282212,0.00585392119111927,-0.0155253298670827,-0.00987485104181107
"3208",-0.0118947214788299,-0.0108620648461809,-0.00440603555050811,-0.00709559586841457,0.00301041347330355,0.00276932722716094,-0.0105836806216673,-0.00657901847039488,0.00547281650006548,-0.000664871068921102
"3209",-0.017664732290289,-0.0261681867118397,-0.012391625894172,-0.00763931480541102,0.00244328396682358,0.00346331171371084,-0.00388975154195093,-0.00560356395196959,0.0116736370524373,-0.0086494124123877
"3210",0.00819283290342265,0.00695780357436315,0.00501882383157293,0.0129128204795237,0.0091218771644741,0.00522123031284583,0.00976235197853925,0.00768440199371345,0.0045306457783747,-0.00134230457842133
"3211",0.0135321022713335,0.00905397540397157,0.0115926782138889,0.00441293463921966,0.00738336363006042,0.00193678747828163,0.00537113172993231,0.0119471118727161,0,0.00806451612903225
"3212",-0.00431471912770232,0.000236196577638292,-0.00634695619869641,-0.00829874887677129,-0.00828830626667842,-0.00333884440071008,-0.00277795189328323,-0.00326547960432411,-0.00852707576576783,-0.0013333559115386
"3213",-0.0155246724927783,-0.0110954095815514,-0.00585524631585277,-0.00713760938652341,0.00269390323263363,0.00211573436804202,-0.00514309522442802,-0.00302420550853988,0.00874259707523506,-0.000667466324014487
"3214",0.00949640708822885,0.00811644237714471,0.00874531607352669,0.00768468867866967,-0.00564855402328646,-0.00255123372670574,0.00323100453966663,0.00505556896077586,0.000916044263191251,0.00267198788324197
"3215",0.00676346735717548,0.00899842411551632,-0.00123852281482706,0.0103320246432104,-0.0148946308303881,-0.00626206512166205,0.00193243515201091,0.00100607596912972,-0.00872935567625432,0.00666220231940717
"3216",0.0103668977558902,0.021121742548367,0.01240040729624,0.0160701558228009,-0.0123766223909908,-0.00683415672789955,-0.000750086793809945,0.0100502465494383,-0.00553937228235746,0.0119126403683329
"3217",-0.00111375540308856,-0.00436681707647868,-0.00437444383659746,-0.00431343189990863,0.00726287291355443,0.00277034766623263,0.000214471384670345,-0.00124377720588753,0.00399912164535543,-0.0045781334059144
"3218",0.00990037166970725,0.0129271410544696,0.0149384778245647,0.00890486456055917,-0.0120883401179357,-0.00481243362713624,0.000536063491396677,0.00697385807325257,-0.00697058843361797,-0.0026280985247561
"3219",-0.00160602718556602,0.000911522426665812,-0.00207797090455231,0.00286263656985342,0.00121643995403198,0.00197001559850785,0.000750000229935432,0.00692545482035012,0.00573026999691795,0.00131747834751383
"3220",0.00294908642414593,0.00478146696455273,-0.00260280208727059,0.00380592940259072,-0.00242991684560956,-0.000357433780777905,0.00556737840711174,0.00147394998266259,0.00142437856493483,0.00394743517647012
"3221",-0.00437716540730426,0.000679757534593373,-0.0019137248191381,-0.00521332050936663,0,0.000894097512452063,0.00798554638770121,-0.000245366442058303,-0.00106673777777744,-0.000655352323614466
"3222",0.00677915091704806,0.00407609380126428,0.00714660775444353,0.0090519864372629,-0.00752266053743211,-0.00366227420716436,0.00728853671727125,0.00588822775426934,-0.00477014072767334,-0.00131149755965509
"3223",-0.00326672069010003,-0.0040595467080915,0.00121149703063694,0.000708128977800593,0.00584711696354767,0.00233092994426598,-0.00325084489201311,-0.000731762150698922,0.00293299964611915,0.00131321984427624
"3224",0.00290953245626957,0.00634054223440583,0.00414868798958046,0.000236028559744694,0.00100471967528759,0.000357649429707063,0.00136765129010241,0.000244064676203193,0.00235379462953911,0.0124589936319914
"3225",0.00163401144780484,0.00360039390117328,0.000516399885898799,0,-0.00200730679798589,-0.00017872927035989,-0.00126078514379435,-0.00390436787364301,0.00711591835989411,0.00518143477574506
"3226",0.00409500551708786,-0.000672616778097268,-0.000516133354693249,0.00707545215445449,-0.00488519485352168,-0.00214619719676801,-0.0102041233680787,-0.00367471017080689,0.00233167527966982,0.00579890297429775
"3227",0.00563649510849085,0.00426287134459868,0.00292641118715453,0.00585476494555115,-0.00909634089728306,-0.00376420747378869,-0.00542026138688778,0.00122950845432102,-0.00860004223459732,-0.00384362468784738
"3228",-0.000296766805028659,-0.00134040244323375,0.00429115214121811,-0.00512228470529752,0.000656017412822063,0.000899583983169583,0.00341954883089657,-0.00122799861963618,-0.00277303045202659,-0.00192926024006812
"3229",0.00306726754808562,0.00626394495282478,0.00273454742982326,0.00444654076114004,0.014634007156876,0.00485353408977796,0.00553772242219464,0.00442596330482825,0.00549022459893056,-0.00644334190948614
"3230",-0.00266332612602393,-0.00333478382964869,0.000170477625216936,-0.00792161431926885,0.0134903371240434,0.00635062577167145,-0.00169443531309976,0.00342722965155584,0.00999850347472697,-0.0058365754909161
"3231",0.00926398060928735,0.00736111691808872,0.00988411997916749,0.0150304810680795,-0.00307817484639594,-0.00188709452282398,-0.000742686186689379,0.00390331107524844,0.000912764209712646,0.0182648168799422
"3232",0.00401772581492499,0.00465017786621624,0.00674989804278514,0.00994914535714386,-0.0131615449648247,-0.0050834062749322,-0.00775030130625542,-0.00121508893840683,-0.0028760101413583,0.00640612793002915
"3233",-0.00110619606818874,-0.00264493869093796,0.00134096918594984,0.00572734148166232,-0.0112466351621066,-0.00537836659918323,-0.0162636261385525,-0.003649571950746,-0.0161800077177632,0.00254619201042838
"3234",0.000228034848657854,0.0013259764719431,-0.00217609112971717,-0.00318918141218405,0.0060517681253045,0.00288395150539,0.00293665833290269,-0.00293038850569194,0.00429024650882015,-0.0107936716004128
"3235",0.00351673976531486,-0.000220766378140391,0.00587145504308784,0.00731274290725459,-0.0181185409809774,-0.00799782172619234,-0.00954339832380979,-0.00269412548072823,-0.0155214884055853,-0.000641891971205011
"3236",0.00246610843398765,0.00022081512669625,-0.000500294710443328,-0.00907444700083282,-0.00420723215131547,-0.0013588085953703,-0.00186135389775088,-0.00982317808616628,-0.00636439556333568,0.00256908653475652
"3237",-0.00190980324376389,-0.00154489809833214,-0.0025029282751281,-0.00709707762687761,0.000667080177745083,0.00108859528762872,0.00230364905490199,-0.00471227623206194,-0.00240192883326229,-0.00640612793002915
"3238",0.00210799455353805,0.00110522832340321,0.00217465200582745,-0.00645605031905561,0.00459258814699193,0.000453031960672368,-0.00700450617708126,-0.00523314608433978,0.00269951120238598,0.000644788954934805
"3239",0.000323648170976965,-0.00198724132789829,-0.00350525584842576,-0.0076584514720679,0.00648874478361572,0.00271712480323383,0.00815608582143668,-0.0055109200775979,0.00400205943399845,0.00193298947981591
"3240",0.00145579275335095,-0.000221214563494887,-0.00435518301594739,0.000701600342905895,0.0103297300349896,0.00505825698692797,0.0079806797187405,0.00428212400562367,0.00420352237146027,-0.00321552085191401
"3241",0.00723638944472116,0.0046470906042555,0.00588838418716042,0.00794580023319202,-0.00108786789634852,-0.000808830076967415,0.00531460881761636,0.00777522933635288,-0.00252591660689849,0.00516131205968251
"3242",0.00073760270939327,0.00132150672653375,0.000836217831834185,-0.00162297612260753,0.00181479306136789,0.0017089475494716,0.00517851987483331,0.0074663781958153,0.00296641327859848,-0.0102695541958202
"3243",-0.000288376463890461,-0.00131976265131262,-0.00317511822330563,0.0020901367221573,0.00833287595610011,0.00188565378545369,0.00128798462890245,0.0037055748916679,0.000505028152684606,-0.00907920528324691
"3244",-0.00371889012992432,-0.00594719046175507,-0.0030175718647133,-0.00440335468351993,0.0103476996316423,0.00367444608778555,-0.000214402409897674,-0.000738426047292018,0.000504672283442753,0.0130890276901821
"3245",-0.00160882372462834,-0.00177270680161112,0.00100883365842619,-0.00209493087638679,-0.0062589160279064,-0.00250022603355515,-0.0137236357518661,-0.00492596221107222,-0.00547704689669382,0.00904394952668475
"3246",0.0022238397447345,0.00244175296572791,0.000671991283627715,0,0.00128833152401819,-0.000179012059175587,-0.00326113395856065,-0.00371291217138692,-0.00188402173913049,-0.000640183169661301
"3247",0.00775024116332945,0.00819308030315824,0.00688260565951326,0.0100303013228731,0.00293078590594553,0.000447637280721169,0.00392622397437226,0.00546586892975909,-0.00479165802266368,0
"3248",0.002265646260867,0.00109827715633704,-0.00166713796179052,-0.00300232900928166,0.00584420628485072,0.00187934693454328,0.0120587404793282,0.0042005448762279,0.00481472855537302,0.00576553466334007
"3249",0.00445748704343796,0.00153574657871358,0.00200397055985202,0.00115829935875245,-0.00290523553139865,-0.00259039765954372,0.00322017687568765,0.00196855552877606,-0.00529991268694952,-0.00509556275296941
"3250",-0.00370863507333941,-0.00569556505851587,-0.0095000378293375,-0.0157334689917172,-0.00213185300371277,-0.000806077040950703,-0.00278197784998413,-0.00294704497579279,0.00620397073950696,-0.0198463287199427
"3251",-0.00849474665826089,-0.00793127564336493,-0.00201914464399422,-0.000235100245813191,-0.013333034970482,-0.00359027587681104,-0.014806828672505,-0.00270925691681523,-0.000507819523372866,-0.00130635779152333
"3252",-0.00670655019481359,-0.00421941390456804,0.00387790695224277,-0.0051727732738055,0.0209675315711753,0.00891808522589677,0.00609883853717097,-0.00197587445505409,0.00957985388677685,0.000654066522213448
"3253",0.00617028188067215,0.00958965082967977,0.0112529604153286,0.0075632594891859,-0.00998520311141649,-0.00383931237076141,0.00389699724798431,0.00222723318939066,-0.00136584716148491,0.0156862734681336
"3254",0.00179795397109284,-0.00176713571407061,-0.00398605851785527,0.00445687497936542,-0.00486419732270682,-0.00233028087990439,0.000862608653534158,0.000987667009547,0.000575885409960897,0.00193043642338497
"3255",0.00913403841683103,0.00885147598331959,0.0115057535348513,0.00583835770721075,-0.00553463755845196,-0.00305455024045198,0.00172380656187587,0.00666014143844662,-0.00992809352517998,0.00642265108196249
"3256",-0.0031440959318807,-0.004386907386289,-0.00560500436201128,-0.00394700107289137,0.00216819498851106,0.000811029707273203,0.00204343999727863,-0.000980190551486126,-0.00029060457384833,-0.00127634574400448
"3257",-0.00111510577620166,0.00044059931886431,-0.000497375950976875,0.00349648210265263,0.0000722054534727512,-0.00117059928357277,-0.00601046847909958,-0.00171693809327855,0.00283470703830924,0.00447288663458867
"3258",0.00283866081989625,0.00484476839009584,0.00215625641740491,0.0146341662473077,0.00786108737547142,0.00414680720751703,-0.00971824170688707,-0.00196565331534515,0.00688553303699702,-0.00445296900902392
"3259",0.00861906234635379,0.00832784148115495,0.0024826298230145,0.0173991890283409,-0.0164579754579107,-0.00790014170982722,-0.0130847032369468,-0.00467747370951554,-0.00352724594770004,0.00894570834782171
"3260",0.000599077641106893,0.0091284730523935,0.00264152806361473,-0.000450028496518762,0.011567723735441,0.00588177194240602,0.000994355607379482,-0.00296807841061297,0.00447887041358164,0.00506645466891054
"3261",0.00687006067188367,0.0133553244871363,0.00459901053747536,0.00848460659570516,-0.00899021143348189,-0.00467796822214595,0.00642044741357362,0.00620188901389418,-0.0000719884917945723,0.00693133829067927
"3262",0.000219137850890005,-0.00706037624902112,-0.00215626136745295,0.00911985843319996,-0.00137879623338311,0.0000904870448859008,-0.00852812040615658,-0.00665683130481187,-0.000215750873923115,0.0043804543080963
"3263",0.0000624735597016812,-0.00107733247145014,-0.0039893949468085,0.00542254882162441,-0.00821233403371502,-0.00271136247232229,0.0129580321590046,-0.000992735676776713,0.000072002016833439,0.000623031858375089
"3264",0.00409899620974241,0.000215660047117039,-0.00100128508014974,0.000449438202247299,0.0015999655557859,0.000780468400041423,0.00827084252315835,0.00844711485816307,0.00258956257834675,0.00435869731147753
"3265",0.00438425471141235,0.00345050686759762,-0.000668242554823784,0.00202158580413281,0.00131901930231626,0,0.00623427758941264,0.00098550337032921,0.00100444106025099,-0.00123988358548832
"3266",0.00152773355531122,0.0023640662446609,-0.000835840855900938,0.00134492263293162,-0.00146368231376826,-0.000906713656492752,-0.00565214130434788,-0.000157316625596371,0.00308194515246707,0.000252270433905188
"3267",0.0000311624430882063,0,-0.0040154090680945,-0.00223859423499417,0.00285830028917866,0.00172440949252328,0.00273283768912869,0.00262199797121121,0.00943199019861352,0.00441361916771754
"3268",0.00532326040981279,0.00385936972254219,0.00268772052221955,0.00717969486201486,0.00241155460169074,0.00144964601975373,0.00534174189441594,0.00679911052305915,0.00785730139853325,0.00753289391086009
"3269",-0.000247776675247557,0.00384451089278093,-0.00184280452073726,0.00400982410358264,0.00109357461654302,0.00144761108026614,0.00271090866719903,0.00649350649350655,-0.000351193975586694,0.0018692213002629
"3270",-0.00551321960818396,-0.0068085106382979,-0.00889565260504688,-0.00665631240292874,-0.00364108166163768,-0.000632409262915412,0.000757002262820494,-0.00206456774193553,0.00210779874787059,-0.00186573383084565
"3271",0.00242929497813882,0.00599826478149112,0.00321766305195026,0.00223361626088892,-0.00979397105818702,-0.00361591550949691,0.00583532520169294,0.00310325850029769,0.00189293269673496,-0.0062304676779108
"3272",0.00935192363225901,0.00787911004853292,0.0104658841841363,0.0202808116844397,0.0112931652637001,0.00462708482368202,-0.0110657389113505,0.00206233560035241,0.00734781696351927,0.00125391849529799
"3273",-0.00757223208625346,-0.0107754485199473,-0.0110257265114312,-0.0185670384134345,0.0154003276662347,0.0066828872442124,0.00716997260717078,-0.00205809112575495,0.0132685240695074,0.0118973074514714
"3274",0.00381505221531531,0.00363096967108056,0.00354728034548502,-0.00244825283774763,-0.00567850982108675,-0.00107653251572137,0.000862927417354387,0.00232018555503521,0.0104894967058171,0.00185649752475237
"3275",-0.0028117783890228,-0.00574592442026267,0.00168318464904904,-0.000669321731370021,-0.00491578757226407,-0.00143688756856275,-0.0101304342048666,-0.00360079723248985,0.00393515166520908,-0.000617726953815456
"3276",0.00532953534339886,0.00192636982178129,0.000168072598490054,0.00580482237542257,-0.0066109623040328,-0.00233831119270489,0.0023952314076261,-0.00722774872339949,-0.00750152052779929,-0.0148331273176762
"3277",0.00678065008054296,0.00299081386475519,0.00705643481182783,0.00665924543083785,0.00351033169113135,0.000721154860710671,0.00054309764309779,-0.000780005220489044,-0.00565165459858608,-0.00439146800501888
"3278",-0.00287770707872714,-0.00489882843665956,-0.00700699044055697,0.00529221633041765,0.00889076978754466,0.00216200485536233,0.00868427023390361,0.00052045277127255,0.00602619328922938,0
"3279",0.00687734813759522,0.00449484151338098,0.00571238239247296,0.01557356876508,-0.00303370324154906,-0.00116859708026729,0.010654391103194,0.00546161234170039,-0.00741948791996483,-0.00756143667296783
"3280",-0.00152462260010533,0.000639228638397604,0.000334112924588847,-0.00561550768068053,0.0051440858471965,0.00197985491042485,-0.00383346805096496,-0.000775969994826653,-0.000891544326973026,0.00444444444444447
"3281",0.00225985638381943,-0.000638820286176012,-0.00367403133476907,-0.00781930912642681,0.00663165376038166,0.00251480604224463,0.00887219640174686,0.00336518241353412,0.00583424386252673,-0.0050568900126422
"3282",0.0083183856405229,0.00554014489665455,0.000670482735501299,0.00634853327495621,-0.00315078069797303,-0.00206055196774468,0.00741687881172526,0.00644994873322746,-0.00156950328228833,-0.00127064803049548
"3283",0.0031125316074494,0.00487389287717499,0.000670033489614141,0.00565584064268343,-0.00854816137614078,-0.000807927497977534,0.00115692046367455,0.00410151264298952,0.00184542412474098,0.00318066157760799
"3284",-0.0019581984530852,-0.00801343348854644,-0.0053566118059386,-0.0253082197707116,0.0105056472041953,0.00395317064646505,0.0101901668202506,-0.0066376822383295,0.00109157455189557,-0.00570703868103994
"3285",0.000120760644277462,0.000637733829980336,0.00454394158680382,0.00821125148221813,0.00351339429654574,0.00017907378827009,-0.00571966490350817,0.00411205345669496,0.000340656932647843,-0.0133928571428571
"3286",0.00114687331619345,-0.00403652007648181,0.00117270901612843,-0.0103456086286594,0.00700187178587486,0.00250535521707218,0.00596170896389814,0.00204765804965445,0.00224812327635981,-0.0084033613445379
"3287",-0.00889307847313081,-0.00234643766325848,-0.00384871164152323,-0.0080071398578101,0.00808853465307369,0.00357015871420563,-0.00228738823040142,0.00229885045727451,0.00584557523944995,-0.0149934810951761
"3288",-0.0160294101539785,-0.020525956809921,-0.0179741309923421,-0.0345290822658781,0.0155546032497662,0.00675914082289064,-0.00479365365562368,-0.0127420992486188,0.00682530765847567,-0.0185307743216413
"3289",0.0104791808346214,0.0087316741163137,0.0088949881781557,0.00836035744634556,-0.00783136575410537,-0.00335695163242944,0.00429323560209416,0.00129062977332839,-0.00892678002125047,0.00472016183411994
"3290",-0.000826027066014867,0.00129844192379225,-0.00322141403865717,0.00483655019974893,0.00977925393376888,0.00478641538297664,-0.00312796358552969,0.00567148735056766,0.00541787199193089,-0.00469798657718123
"3291",0.00324535550862404,-0.00129675815863406,-0.00136080963835994,-0.0148980285377487,0.000138389818672868,0.000970401833170431,0.0012551197442201,-0.000256293271278851,0.0000673177928653956,-0.00876601483479433
"3292",-0.0181579044406291,-0.0157974251416886,-0.0163515417535607,-0.020241949744067,0.00912982069713131,0.0050233749974995,-0.0121174445173683,-0.00410256410256404,0.0057924226726449,-0.00816326530612244
"3293",0.00742853920456943,0.000879507475813668,0.00761903030303035,0.0111612678422877,-0.000810130567652001,-0.000851737342510206,0.00306652215290271,-0.00102989186405777,-0.00649568731673889,-0.0185185185185185
"3294",0.0152412781568751,0.0158172671353249,0.0151228907909071,0.0258336765695784,-0.013467075134852,-0.00580021085724769,0.0102256060486443,0.00489698466229327,-0.0130089511120994,0.00139762403913335
"3295",0.0115480065127818,0.0114618939679112,0.0089723717623158,0.0057234432234432,-0.0109346916514019,-0.00433125643181542,0.000208661166468671,0.000512849422269923,0.00122931099231849,0.0153524075366365
"3296",0.00336485624728966,0.00171045542014103,0.00755035260236081,0.000910562258138015,0.00450670172773182,0.000710214066304005,0.0037558790559391,-0.000512586542557814,0.0053883977533018,0.00412371134020617
"3297",-0.0053296572889806,-0.00875131307369525,-0.00965858467374825,-0.0138730949767322,0.0124780915111904,0.00479067364842334,-0.000415767596047778,-0.00461659376165191,0.00264585492452607,-0.00547570157426425
"3298",0.00746532483568974,0.00258402245012967,-0.00117704723092238,0.00553498603470981,0.00276963830886379,0.00194240379466293,0.010086316108689,0.00566859042338064,0.00257124986804746,-0.00894700619408118
"3299",0.0017330495163479,0.00601372409764345,0.00505048804543806,0.0130733950951099,-0.00504042226730006,-0.00237925941770123,0.00813260251320358,0.00358695884158244,-0.00344195185856722,0.0034722222222221
"3300",0.00644276959843793,0.00576432536293758,-0.00485763810958739,0.0135839263565283,-0.00506594987903297,-0.00256164861860475,0.00796486265699969,0.000510620398806338,-0.000812752246708404,0.013840830449827
"3301",-0.00106696397999362,-0.00785393742615292,-0.00875275206194237,-0.0131784677239224,0.00383626271841164,0.00088555075130925,0.00678753932517018,0.000255218174412208,0.00569345289314205,0.000682593856655256
"3302",0.0016021123930583,0.000855733810195325,-0.00747152330568057,0.000452716161158939,0.00437745220694152,0.00247747584941616,0.00905616851648738,0.00867346916649314,0.00417842687092507,-0.000682128240109159
"3303",-0.00257699936178324,-0.00448907662439235,-0.0148844993176305,-0.00656110844884383,0.00684874220770793,0.00158871943895322,-0.000698045479637588,-0.00354069287959791,0.0128188187919462,0.00750853242320826
"3304",0.00478123406707587,0.00579772385656008,-0.0017367488108111,0.00728763379640163,-0.0000686734762954666,-0.00017628555164384,-0.0125736155331166,-0.00304576126671274,0.00583121712726231,0.00948509485094862
"3305",-0.00410824619150252,-0.00597777540563627,-0.0064370041753653,-0.0156002486999774,0.00783344979494038,0.00290856705236608,0.0108135425208755,-0.00381868645159578,0.00408466320964895,-0.00402684563758393
"3306",-0.0102982664384058,-0.00279211763762632,-0.00840483263167857,-0.00574184644598419,0.00934060165826422,0.00404252747704481,0.00189964012896326,-0.00204451822017593,0.0150252144865768,-0.00404312668463613
"3307",-0.0331654001294849,-0.043291018737885,-0.033727705567231,-0.0374221058576552,0.0149285049831758,0.00778987821556121,-0.0133718791874252,-0.0197183103641053,0.00898512622466319,-0.0189445196211095
"3308",-0.0303021481486014,-0.0229625404305511,-0.00164473681204802,-0.00791931883462049,0.00532450983399424,0.0027792346298483,-0.0268028918740905,-0.0107105540937971,-0.0178742588986933,-0.0186206896551724
"3309",-0.00367821532726464,0.000921589819281587,0.00494235758846129,0.00798253507498781,-0.00529630958154337,-0.000519605324021732,-0.0104967988931948,-0.0105623979551728,0.00437050219757662,-0.00983836964160234
"3310",-0.0449116853932584,-0.0303867410310024,-0.0342441153280831,-0.0239980813054035,0.0108485684762554,0.00485263940165948,-0.0524104406302955,-0.0240192414192891,0.000194836655226238,-0.0170333569907736
"3311",-0.00420153930282885,-0.00807217493048862,-0.00113166729536018,-0.00368817328193616,0.0225836157201298,0.0112108240860327,-0.0312569160800608,-0.0213289308176101,-0.0364934740259739,-0.0173285198555957
"3312",0.0433065063354314,0.0179511732396165,0.0126510954050434,0.0217177196446199,-0.00735739416269166,-0.00068307716829541,0.0481693238405188,0.00558818090002289,0.00552629715843445,0.0227773695811904
"3313",-0.0286324569365876,-0.00893479917551832,-0.012865970298975,-0.00676335716119048,0.0155255292253407,0.0116199674331854,0.000109180219308058,0.0133370095394829,0.0314343303907707,0.00215517241379315
"3314",0.0420330249811161,0.0360615878499839,0.0217227242486349,0.0177528944006053,-0.0106185887466439,-0.00219597124668969,0.038201264848245,0.0235810522736206,0.00175453246965063,0.000716845878136363
"3315",-0.0332416879710583,-0.0316005739226277,-0.0181179330745056,-0.0210274084123013,0.0248917440342891,0.00888778575324012,-0.0217619841748743,-0.00375041501471118,0.0216009400207333,-0.0107449856733525
"3316",-0.0165311120438405,-0.0151335773200856,-0.00960276765952228,-0.0205028064314668,0.0520439048184733,0.010151858207033,-0.0169801391623814,-0.0188221838887386,0.000380963858627181,-0.0325850832729907
"3317",-0.0780944688457279,-0.087154905778876,-0.0509505722794894,-0.0682781443239934,0.0271031294092912,0.00897010782441687,-0.0741226514253562,-0.0570019700190754,0.00165023798825326,-0.0778443113772455
"3318",0.0517448908974445,0.0360336401893739,0.0298477976701841,0.0508157809792933,-0.0512580907163678,-0.0183569554241779,0.038611369970212,0.00610284800929972,-0.0211013373183111,0.0316558441558441
"3319",-0.048748447979579,-0.0558517404379727,-0.0338455942423652,-0.0465767868013033,-0.0367977120422655,-0.00997905241090158,-0.0582083112574842,-0.0283073376171963,-0.00356035094666884,-0.0180959874114871
"3320",-0.0956771593350247,-0.113471312542923,-0.0980470947472154,-0.100106783238302,0.00619690159200736,0.00050825852123082,-0.0974166995372621,-0.103448249210709,-0.039888262711738,-0.0400641025641025
"3321",0.0854863000867101,0.0606612053181315,0.032812523053851,0.0720854367275419,-0.022603161904762,-0.00651883661059505,0.0853284105387886,-0.0135941644562334,-0.0305162339374359,0.0108514190317195
"3322",-0.109423734717191,-0.113239945289107,-0.0659174194942728,-0.124792477166366,0.0647655051998766,0.0264166941016906,-0.16869997119655,-0.09882356302521,-0.011446119566207,-0.060280759702725
"3323",0.0539920645238592,0.0451467268623023,0.0490513408363873,0.0689219749896293,-0.0666829829373928,-0.0250726199685998,0.0469907804178888,-0.019395673979697,0.013555485834196,-0.0158172231985941
"3324",-0.0506329226586283,-0.0688059240975006,-0.0211733348037054,-0.0863650373745922,-0.056412539061643,-0.0138805841778081,-0.0984000749709787,-0.0928109892426402,-0.0199219910827807,-0.0330357142857142
