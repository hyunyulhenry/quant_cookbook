"","SPY","IEV","EWJ","EEM","TLT","IEF","IYR","RWX","GLD","DBC"
"1",0.00212204857892062,-0.00568168217719622,0.0105634253417877,-0.0138089105329995,0.00606396543910592,0.00362832452924011,-0.000238518041803526,-0.0074364728506715,-0.01011555892928,-0.0260503050587256
"2",-0.00797636883866415,-0.0147620707440701,-0.0257840909953339,-0.029238232118335,-0.00435324775908241,-0.00325396988848048,-0.0155035981684098,-0.0124343117072752,-0.0240065523436642,-0.0034512995305368
"3",0.00462528813875518,0.00164359391516467,0.00572274003685114,0.00725729202176173,0.00179378784542861,0.000725244422058013,-0.000242183735400303,-0.00338955372229766,0.00515210254785115,0.00519471605092869
"4",-0.00085015723037718,-0.00376392258712888,0.00640078219274787,-0.0223362924377141,0,-0.000241179499985478,0.0117532150387523,0.00161926858631745,0.00611769179894184,-0.00861317890472024
"5",0.00333187221950659,-0.00561869664923631,-0.0148409764866628,-0.00230322563786678,-0.00447656887763093,-0.00169193183234639,0.0159282760840618,-0.00565985269618152,-0.00427276924479103,-0.0147698688123383
"6",0.0043803417871402,0.0108136444671405,-0.00502146472722409,0.0126500976777097,-0.0058433058231081,-0.00266323648224698,0.0114346314523921,0.00325279468212258,0.000660191450734482,-0.00132265790941177
"7",0.00759702246868055,0.00905916064364232,0.0129778439592207,0.0203336510059355,-0.0046355940689764,-0.00206330406739019,0.00349637356292964,0.00664595616707353,0.0253999171136414,0.0233996224013486
"8",-0.00195453187590677,0,0.00355863118259458,0.00357479476500355,0.00215861864754952,0.00194630286406094,0.0114982279379352,0.0025765238900326,-0.0032169375331168,-0.0228645994088241
"9",0.000419676336849362,-0.00057320548157358,0,-0.00418510565721741,-0.0030614950425405,-0.00194252212768031,0.00298526677483646,0.00706733772156154,0.0108116506243077,0.00883002834000157
"10",-0.00335606724273252,-0.00305805850170693,-0.000709071161415498,-0.0105519126638738,0.00307089657718773,0.00133760750089307,-0.0034341924237602,-0.00111644408223477,-0.00606642729991103,-0.0105032427762808
"11",0.00196413908577542,0.010736529498701,0.00709712247323369,0.0179848978084849,-0.00272088740150667,-0.00157822034597566,0.00884487158636627,0.00973966460559961,0.0118856733660673,0.0150376039605462
"12",-0.00308047641444475,-0.00701844334953416,0,-0.00115420872356675,0.00238638942762592,0.00182415241669065,-0.00307381089273506,0.0102783903576438,-0.00444442857142857,0.000871366900456527
"13",0.00294969164484793,0.00897803144092069,0.00563765618722312,0.0227531712362872,-0.00657588438954526,-0.00291398629690731,0.00285533512446756,0.00751297955584795,0.0240752866059424,0.0317805604448693
"14",0.00805306455854971,0.00511174160021977,0.0133146661703822,0.00869064961107013,-0.000113741406236545,0.000121291705275084,0.0136675773965071,0.000931827879582681,0.00155688923134556,-0.00843882505047222
"15",-0.0117403214149138,-0.0154452588873589,-0.0165974452142039,-0.0307572440750817,-0.00719195653401017,-0.00389667434478425,0.00595539476785145,-0.00589734210841641,-0.00419717070737846,-0.00893599478055107
"16",-0.000913619243186337,0.00277407153825426,0.000703326089980916,0.00613329097049053,-0.000803958058334664,-0.000121630258104855,0.0030154113562153,-0.00624547015638688,0.00171714023469072,0.0124515654514379
"17",-0.000562882915589369,0.0022893137961153,0.00351370355008207,-0.01325243548375,-0.00218567677253401,-0.000734198096313032,0.00289480662208241,0.00612762787039611,-0.00623341144564171,-0.020356203459988
"18",0.00520934466799239,0.0053297136940591,0.00630247366792824,0.0154895962540875,0.00115242710820085,0.000978985972805102,0.00344265441994107,0.00405983617508987,0.00705662537243201,0.027705554222162
"19",0.00672330041230507,0.00511190979089271,-0.00417528408218704,0.00775912267216516,0.00840761602030282,0.00366730831884965,0.0113977351343699,0,0.00949861399099006,0.0105308029970261
"20",0.00598240425763352,0.0078180500002436,0.0132771437257546,0.0122479853999327,-0.00120360960283983,-0.000721801178719561,-0.000547532375871018,0.0113528300567416,0.00601571784619104,-0.00375161049023653
"21",0.00138307910778601,-0.000934844588558859,-0.00620695784488834,-0.00302487826939379,0.00126275701914014,0.000856419605227421,0.00711554384543511,0.0110719112766913,-0.0144127872675132,0.0129706315284444
"22",0.00027622826730922,-0.00327404071351867,-0.00763325208825449,0.000953722565128823,0.00137546453058346,0.00110032388684211,-0.000651883880573578,0.00304185694023773,0.000466692602157481,-0.00330437818714768
"23",0.00027629864165446,0.00656978941267794,0.00839153072221488,0.00987341364191252,0.00549808930522522,0.00280807317248155,0.0137043662635137,0.0103103523047769,0.00746389387230284,-0.00497302215289619
"24",0.00220850485816459,0.00372958970222959,-0.000693742351985382,-0.00385925540833332,0.00296115530164309,0.0021925715571911,0.0146998441098405,0.00405252116642107,-0.00246957860056218,-0.0120781760068096
"25",-0.00130844241645078,-0.00232225488499993,-0.0124910213879003,-0.00533802395976535,0.000795312466929099,0.000241934119855181,-0.00761369799104561,-0.000598028930855032,0.0137706953630217,0.0231870629732278
"26",-0.00744734420744309,-0.00595933577643581,0.00281078505617094,-0.0119448339366696,-0.00567427558569111,-0.00303632860864977,-0.0141714466608379,0.000598386783463356,0.00915760115190478,0.00618051849681645
"27",-0.00340413788116178,-0.00327833440786018,-0.000700883418384257,-0.00683305353893715,-0.0022811981331391,-0.00133972898503254,-0.0167531476330951,-0.00822136618038116,-0.00680588293379225,-0.0188371198035659
"28",0.00843474458263116,0.00977369880003387,0.0210380696172994,0.015877111670759,-0.00217402617908613,-0.000732306324060517,0.0178080441590702,0.00813881663311311,0.00258867070469515,0.0183639546801622
"29",0.00656734450623131,0.0128431825558735,0.0164835566505572,0.0215334747581035,0.00951397741218152,0.00573849967579387,-0.00615623749305394,0.0165944620333944,0.00804992454738307,-0.0135245569450847
"30",0.00130450162889684,-0.00202139091666986,0.00810820050638994,0.000594712210308046,0.00295253018419039,0.00157755391581071,0.00825918734862241,0.00294123737616503,0.00060269697441484,0
"31",-0.000479661969168377,-0.000276243070824078,-0.000670493556458762,0.00229402859702277,0.003509674434927,0.0010911938819429,-0.0034488161985311,-0.00073359923156846,-0.000752943788408844,0.0174491644849777
"32",0.00212696249666577,0.00349936734538669,-0.00335328933917156,0.00262725484045823,0.00225646493184839,0.00121052979398506,0.00843595564697663,0.001908258082572,-0.015822829779644,-0.0110249158425911
"33",-0.000410825445496532,-0.00734186828056127,0.000672723335915615,0.00295816149657702,-0.00168865924228012,-0.000121283550759466,-0.00525533221647123,0.0032215221571843,0.0312356463400902,0.0214698305811687
"34",-0.000753221233364521,0.00286606170062509,0.00269003873391016,-0.00252838464507532,-0.00541216967768321,-0.00253982629119964,-0.00506728273361867,0.00627739097785063,-0.00296950268654794,0.013742936552138
"35",-0.00390797597636028,0.00258146656705249,0.00871907786281323,-0.00718192631172043,0.00714234087418197,0.0040015259120223,-0.014196052174536,0.00681873641717501,0.00848844352975586,0.00637963267720099
"36",-0.000894358193119893,0.00505730587081632,0.00664924485183693,-0.000425442882123872,0.006641705716671,0.00313944072429018,-0.00648548202463683,-0.00806919656855454,0.00561129643220171,0.00277337747782158
"37",-0.0390580504486641,-0.0539797168578178,-0.023778418053093,-0.0813113014527554,0.0126346670429609,0.0084265670282746,-0.0324191452078957,-0.0368971680434145,-0.0395006472687415,-0.0189648488774585
"38",0.0102511611428888,0.013539775966515,-0.00135320946228379,0.0250232290957992,-0.00452749551430098,-0.00346164011722749,0.00777638634604272,-0.00558101754437623,0.0163583387030521,0.0153039919303792
"39",-0.00298011689334943,-0.0131680518500058,-0.00474249414971772,-0.0143761778923288,-0.000633731023447437,0.000901406407904703,-0.00624101474749172,-0.012133598345716,-0.00992784251228152,-0.00713994426755238
"40",-0.0130953442510479,-0.0130537743108291,-0.0163377482796957,-0.00926540650092744,0.00501307346622681,0.00324230264158554,-0.0206670034463701,-0.018885825341054,-0.0320571406867212,-0.00918906513063011
"41",-0.00951871856001474,-0.0202800837490064,-0.0145328589253809,-0.0256479520714373,0.00166275696216989,0.000598489681807868,-0.0354435076031052,-0.0228478056614959,-0.0122429604809757,-0.0149191936410714
"42",0.0171089449231669,0.0276000909739753,0.0238764931352637,0.0439037151034469,-0.00298850080937196,-0.00131591329673286,0.0344496328366957,0.0281869730822666,0.0193866518353727,0.00941465989397505
"43",-0.00100170713134218,0.00194639301743615,-0.00205764739126746,-0.00609912818573599,0.00388550618561734,0.00179620382019174,-0.0142556286422272,0.0118380434471714,0.00233828519600054,0.0137874316339257
"44",0.00845530334759625,0.0103921255872108,0.00893489215386367,0.0258288661571631,-0.000884610309613287,-0.000119710387593952,0.0160030070495338,0.00369442672213816,0.00279937778540984,0.00160000109706515
"45",0.000283999376097688,0.00288381660390669,0.000681056018906778,0.00178601377968279,-0.0105143205519407,-0.00561875742416817,0.012249961933205,0.0111961544792041,-0.00356704387870443,-0.0131789655455684
"46",0.00149142926128909,0.003834177238623,0.00816900015215993,0.00490167653800033,0.00391570702122013,0.00276466368414696,0.00507179948484549,0.00712903990622649,0.00186775097276271,-0.00930789262729326
"47",-0.0194335729675158,-0.0244439267884355,-0.0182311416261993,-0.0290906787890729,0.00601572895721358,0.00443743802447916,-0.0263758728770129,-0.0191262861944046,-0.0100979022791097,-0.00776139923920816
"48",0.0074502312824416,0.00371947589208732,-0.00894097357970436,0.00822137586716831,-0.00454104340011552,-0.00131333258407573,0.00471118785896851,-0.0196534118862111,0.00345257370601737,0.00205841743606472
"49",0.00136363604733014,0.00477795658683089,0.000694223964551322,0.00815433600591664,-0.000110656703998568,-0.00107553318555587,0.00750273496653686,0.0117463042588273,0.000625602136778314,-0.00616274323701982
"50",-0.00279960020235481,0.00349384623222027,-0.000693742351985382,-0.00853789356982582,-0.000223171348384232,-0.000119959501134081,-0.00558520836514864,-0.00346399559345412,0.0100031728665209,0.00248040983341546
"51",0.012055257349447,0.0149902937247959,0.0111035583254859,0.0219364008281735,-0.0021140297456721,-0.00131715517635356,0.0100631227372558,0.0194856548840034,0.001856932751922,0.00494845688755019
"52",0.00549176233291915,0.00981412993687214,0.00892247888166886,0.00656381508983217,0.000556750796971706,0.00143902448804933,0.00324441443030832,0.0151371857308402,0.00818657733044725,0.00123089067396864
"53",0.0164576774644116,0.0245330683655272,0.0108844225014104,0.02996082428449,0.000447309243236882,0.00143577894919722,0.0140867265550426,0.0227445661451007,0.00842658227791837,0.00163947728165459
"54",-0.00076792911960788,-0.00653896440919111,0.00134592419287061,-0.00427777817565023,-0.00791176998858989,-0.00334638933219789,-0.00079634923002958,-0.00589086577830722,-0.000911546642357819,0.0163664913648924
"55",0.00146676931077794,0.00519128514721312,0.00134411511581822,0.00463996320726201,-0.00280800506334999,-0.00155917919022142,-0.000264366462635168,-0.000444485447961607,-0.00927615543564009,0.000402619932218462
"56",-0.00132501694879739,0.000737610626238672,-0.00536932640600118,-0.000598493306080194,0.00123897110808047,0.000841122339488409,-0.0155084927493504,-0.00340888750680213,0.0105908515551543,0.00442656260043939
"57",-0.00237440529048438,-0.00608216940733575,-0.00404858805291286,-0.00445035876103195,-0.00168647150894563,-0.000240282569873074,-0.00828464370020887,-0.00654346572507636,-0.00212635189102994,0.0028045321486756
"58",-0.00727978242752347,-0.00917953194848287,-0.00745249677882798,-0.0178804322249435,-0.00202881770703556,-0.000119140901132075,-0.011648452992868,-0.00748472984536486,0.00532733662073093,0.00958850037405323
"59",0.00105747015139346,0.0103872763881305,0.00136504892255407,0.0198690239044343,-0.00135435886253432,-0.00144216311811385,0.00535746177948915,0.00829491269040239,-0.00605603303303415,0.0193905524746216
"60",0.00021156124448396,0.00342706367868484,-0.00681652937974364,-0.00017142459284103,-0.00192264987984236,-0.00120101182559296,0.00935398709545843,0.0127148980181369,0.00137084535046927,-0.0147516879941152
"61",0.00112661031740058,0.0035998589942996,-0.00549085396576809,0.00686667247828132,0.00165962105558304,0.0011119689259167,0.0118497314257584,0.00531777099806963,0.00167325834113963,-0.00985019969883938
"62",0.0107629039216937,0.0129681226327318,0.00828158451963668,0.0163682654263222,-0.00124796322381038,-0.00084445854438675,0.0086954014023064,0.00573038101891399,-0.000303659842176507,-0.00397922538928086
"63",0.00111342393759783,0.00254191215515709,0.00752932836972731,0.00629073986121909,0.00102237277861916,0.00156994150998635,-0.00655182551581956,-0.000876957972832493,0.0148867684980474,0.0111865837697289
"64",0.00271121613886027,0.00443782841535456,-0.00271736630133368,0.000917061412891051,-0.00374584370151909,-0.00253348460718528,0.000809576117464461,0.00438692379958261,0.000748435885299825,0.00197546276217331
"65",0.00138653027871127,-0.000991931894221532,-0.00136242728314706,0.00574639468137783,-0.00660963770847089,-0.00459403550177873,-0.000693719139699955,0.000145526353868997,-0.00493571634855339,-0.0102523310478511
"66",0.00117672205651798,0.0072203537070068,0.00341064140152136,0.0047195679481693,0.00298236368456117,0.00206511015553779,0.00254535581825288,0.00611395457059905,0.00946948759160504,0.0139442326305543
"67",-0.00408000586883039,-0.00394262629305087,-0.00407894624799499,-0.00923021413429825,-0.000686474822177763,-0.00121289727741369,-0.0133855843470012,-0.0111404952092401,-0.00119121493798613,-0.00157179448515576
"68",0.00444377711109945,0.00710680048118517,-0.00136521739771356,0.0167194063552802,0.00022902272572134,0.000971370381223524,-0.00526276101475076,0.00555969941190781,-0.00134174116452757,0.00590315003881492
"69",0.00456250496967803,0.0074140756705634,-0.00820224952729787,0.00490882206640553,-0.00308913338051431,-0.00169727649808071,0.0109349092364661,-0.00334627609187088,0.0126884314879365,0.00547739648670853
"70",0.00949596077201131,0.0117040718340264,0.0144728256496867,0.0118862419501986,0.00550913969090772,0.00109322378305121,-0.000233108772890844,0.0157660463727354,0.00825480591125038,-0.00778202330855171
"71",0.00265895145255479,0.00131470434447545,-0.00611425233159557,-0.00539091421348437,0.00559418982320925,0.00424567884251692,0.0143092744704094,-0.00546109897937164,-0.00584798228514671,-0.0101961268708496
"72",0.00122377964716236,-0.000525185967262032,0.00136708376425276,-0.00744197339616703,0.00499462285845254,0.00229529470422118,-0.00355585223079635,-0.00173405956055872,0.00558819117647058,0.000396154335922549
"73",-0.000271977820230251,0,-0.0047781871841156,-0.0080682011694857,-0.00169440784630026,-0.000120411962845846,-0.00863235206712609,-0.00376390423506989,-0.0124305065412623,-0.00277227922738532
"74",0.00944102783847778,0.0079690685551661,0.00411516781951216,0.0119131888140394,-0.00260288813072629,-0.00108388881460475,0.0109139566430321,0.00624842802153558,0.0173256036920717,0.0138999306258629
"75",-0.00376789797586496,-0.0056472491049715,-0.0109288842477866,-0.00397844786225587,0.0036307673302467,0.00205055281377553,0.00849882403583457,-0.00216629379295341,-0.00640458543251454,0.00665883749617335
"76",0.000405191622500523,0.000174967691151107,-0.00138124551668362,-0.000163089029761254,0.00372984382770514,0.00192714240431036,-0.00683333901902516,-0.00723592452552824,-0.0077644152427655,-0.0136186866940441
"77",0.0091815223031011,0.0105700608471637,0.00553247462603146,0.0123930360266571,-0.00349109425107164,-0.000601691168437113,0.00137624201142672,0.00918416853502046,0.00236226181770594,0.019723922310988
"78",0.00113765778650765,-0.0031115878620962,-0.00481425123780976,-0.00265777461695527,-0.00723277338782158,-0.00288625894376981,0.00137373485066239,-0.00548934738281359,-0.0150242453236743,-0.00696329557888986
"79",-0.000802232522035706,0.000259670828636427,-0.00552862975224955,-0.00500655386757631,-0.000226923604053408,0,-0.00331541726947771,-0.000726146419039786,0.0103184532532472,0.00506419748851039
"80",-0.00829246790529869,-0.00390087463939415,-0.00764411673989895,-0.0193146938187584,0.0104745335657161,0.00434185275873866,-0.0191603176060033,-0.002180139824003,-0.00695680896852591,-0.00891469419041446
"81",0.00256267349553996,0.000261120647830015,0,0.00397193451237388,0.000723843851143213,0.0000485025330632105,-0.0052639424567712,-0.00335029292605882,-0.0059620513317663,0.00195550177609105
"82",0.00585203890527319,0.00539444368849584,0.00560201637329993,0.0198647814677515,-0.00056571063440658,-0.00120560955376869,0.00823120786177611,0.0201694784778645,-0.000449812552112516,-0.00780644828912236
"83",0.00541668663435213,-0.000865278962998262,0.00139287403059196,0.00840541200597533,-0.0022605614952681,-0.00108592055301182,0.0039653661696859,0.00286537159367262,0.0124511543683676,0.00472082218868608
"84",0.00379110763408574,0.0121263892657799,0.00347705193779824,-0.000320433851792035,0.00407939001480884,0.00253767598644083,-0.00499532963620131,0.00628566769156058,0.0103719665245805,-0.00195784038455937
"85",0.000198682002445105,0,0.00485086440371241,0.00649428449086176,0.00270861820711965,0.000843403362231099,0.00093406381877692,0.0052528563014298,0.000879865057050289,-0.00470760579377849
"86",-0.00132495815378686,-0.00898592994899527,-0.00206885119235711,-0.0129839838676415,-0.00225103052759201,0,-0.00653210231199708,-0.0121453051920888,-0.00542128937728936,-0.00630683405612698
"87",0.0027193655778619,0.00276370957584571,0.0124395448707471,0.0161405378958419,-0.00394862660900652,-0.00325191935409341,0.0116240789324666,0.00114352895486602,-0.00633470858874685,-0.00515664530307158
"88",-0.0104519555789591,-0.0201517759199789,-0.0150170544245314,-0.0244616975307825,0.00237864351793049,0.0025377078161819,-0.00998154043531263,-0.00756828701949352,-0.0214973619643007,-0.00398732915969924
"89",0.00855707109248227,0.0168746010280143,0.00762292742032855,0.0254006357902286,-0.00350266686015555,-0.00204839111132504,0.0111374440638834,0.0141007231080379,0.00681813636363637,0.0148119473263204
"90",-0.00218749363092841,-0.00216068057945307,-0.00275109164468201,-0.00992467184964263,-0.00260779986577264,-0.00144932802251663,-0.0104350970699947,-0.00397277154726183,-0.00255828453987728,-0.00355029840873888
"91",0.000265622081511818,0.00259816362035492,-0.00827572392823128,0.00120308097148203,-0.000340896427955095,-0.000120147099727852,-0.0134741955569317,0.00284916056142892,0.00392278219557607,0.00989703519012286
"92",0.0068409538502594,0.00216024475939269,0.0020860294874876,0.0144975042164637,-0.000682387054298128,-0.000605126885487639,-0.00926372419148624,-0.00724444091890808,-0.0141268858712521,-0.00980004381165411
"93",-0.00197928646678391,-0.00172431394883688,-0.00832732618178811,-0.0036318182293692,-0.00409742838505878,-0.00266261055156702,-0.0179813332477217,-0.00887118914632656,-0.00823170756803993,0.00831350277362031
"94",0.00872494150675407,0.0125217061781457,-0.00279922101798868,0.00515054596944098,-0.00662781678622337,-0.00291176053881215,-0.00866660224219185,-0.00389730532460486,0.00707038140394678,-0.00157051832110122
"95",-0.000524705578692664,-0.00759061142479722,0,0.00181348639420809,0.00299060412178909,0.00133906320715504,0.00689543105019608,-0.00130481947198891,0.00228939265671824,0.00983104263365253
"96",-0.000786244825754956,0.00120292647415643,0.00982462372666704,0.000157304499523558,-0.00516067504611673,-0.00279534154387961,0.0103954744686452,0.000580921952685332,-0.00715701255236845,-0.014408109306017
"97",0.000131333348349028,0.00472108463312138,0.00138962695736078,-0.00157376517442231,-0.00288205787585538,-0.0019503180719449,-0.0078676488603181,0.00203027227571084,0.00521478551601784,0.00474108523167938
"98",-0.00905302941875408,-0.0105936111274619,-0.00485751237790077,-0.024034896052214,0.000924939614604048,0.00134355648217954,-0.0152495911369567,-0.0123029817097307,-0.0120537227333885,-0.00550522883832627
"99",0.00417062684144454,0.00682165819689384,-0.00418401913082955,0.0153414235251754,-0.0023107895422112,-0.00109692010420459,0.00631816501127824,0.00029329796809896,0.00293439382239402,0.0122577335130811
"100",0.00362546082071979,0.000428535689447118,0.0105040939731484,-0.00341972649570177,-0.00011590527799854,-0.00207565656546393,0.0305305251119892,-0.000586098115259337,0.00200181700025182,-0.0218748918446232
"101",0.00814518421797694,0.0048866553702398,0.00207895105036227,0.0102137877001243,0.0020845902519866,0.000978404666401866,0.0255643327304997,0.00630326419324367,-0.00537880743814345,0.00958467109811956
"102",-0.00104214410458725,0.00153545712582792,0.0096820066184613,0.00284384744350641,-0.00184914363420019,-0.000365910170434192,-0.00267876113353849,0.018062406561407,0.012669962721416,0.00909802267606286
"103",0.00495713629458261,0.0089435484338849,0.00547948621258487,0.0249686632458581,-0.00525274220599525,-0.00430887232455823,-0.000467084056188227,0.00300471002029967,0.0137320870654245,0.00744810721222477
"104",0.000129454907893622,0.00303958879501076,0.00340559533986684,-0.0044568614860373,0.00455676299671692,0.00160345287506836,0.00630965560795516,0.00699056402063847,0.00150510230267598,0.00894950605841682
"105",-0.00395858648526848,-0.00547108354309545,-0.00135740519956895,-0.00347405912952825,-0.00628111004111209,-0.00320066024038879,-0.0173013323029705,-0.00878355773901729,-0.00255482412752006,-0.00385662185426483
"106",-0.0107500671991745,-0.0198038671745782,-0.00407894624799499,-0.0251741202996553,-0.000467486983876664,0.00049399432231656,-0.00626244983430291,-0.0195799319777034,0.00060269697441484,-0.00038718847866448
"107",-0.0180454489670464,-0.0231390174051522,-0.00409556795556132,-0.0154151092967592,-0.0179159502051867,-0.00999640091909293,-0.0309158288519026,-0.0236151323284872,-0.0173166982492577,0.00503486046064849
"108",0.013011938736573,0.0142300399646869,0.00479790048980067,0.0176739464647513,-0.000834553966087337,0.00186969263760695,0.0164414314998811,0.00104487271594467,-0.0159362698150086,-0.0177263688049796
"109",0.00172096286890144,0.000435866729777024,-0.00136443333884284,0.00856448822043898,-0.00286444045750911,-0.00261272972683724,-0.0147268085769289,-0.00372796120775742,0.00747424466717161,0.0192232805596453
"110",-0.0109052088682637,-0.0164634527734434,-0.0129781830724933,-0.0173767698251375,-0.0144805310817089,-0.0071105346846535,-0.0210729099912581,-0.0176644394547724,-0.00927355529861917,-0.00269446454548161
"111",0.01496831459017,0.0172704538792645,0.00276814123724867,0.0200052187941349,0.0119005149833402,0.00326635238043305,0.0215265367628859,0.0118865398930532,0.00670828414066427,0.0127363633446651
"112",0.00638619580796029,0.0094897729915786,0.0013804628113625,0.0156894159899599,-0.00252032135590818,0.000250584418549415,-0.0102914251122903,0.00135499807753425,0.00108475129528518,0.00952748724430674
"113",0.00568984765726266,0.0125053227610008,0.00895920322116273,0.0227853091506449,0.00685773180249294,0.00438212803660076,0.0151026759725863,0.00811284466027429,0.00386996916006099,0.00604001949708444
"114",-0.00117604179434949,0.00212928982200911,-0.00204923560336179,0.000905916094356085,-0.00203090190986033,-0.000498216334251955,-0.0148779786814335,-0.00330946061417603,0.00154200467361609,0
"115",0.00248561691598548,0.00144532021519517,-0.000684234832046604,0.00113209602837028,0.00933849590281888,0.00486337097573775,0.000990289774905451,0.00739523711683621,0.00816021592733862,-0.00975602421892541
"116",-0.0138975281432263,-0.0129861537535383,-0.00684952681784645,-0.00851647264986632,-0.00806666931514333,-0.00322641741183727,-0.0178083320762902,-0.0112362440008836,-0.011759376370218,0.00113671378480618
"117",0.0055575506599701,0.00610553760804522,0.00482768116214305,0.012466122307734,-0.00478282632068083,-0.00124631601181369,-0.00402962324000056,0.0037880988384007,-0.00231804979629191,-0.00454197639049791
"118",-0.00940879151458618,-0.00965822393561055,-0.00960874033976722,-0.0132131533608085,0.00648851829676733,0.00299348433222835,-0.00379273978220651,-0.00981144665042721,0.00340769837074673,-0.00228145187285711
"119",-0.00478198276228592,-0.0027617525294793,-0.00554397636996629,-0.00760810205296658,0.00549278183229673,0.00323110652975833,-0.0227155168001898,-0.0213410321894127,-0.00540288677682743,-0.0038110602241177
"120",-0.0102786743742347,-0.00519251212505289,0.00139375847234424,-0.00873992677758118,0.000235938072095321,0.000247983216749237,-0.00142836112183742,0.00233659557967791,-0.0125717988514669,-0.0114765510385546
"121",0.0142290923362984,0.00913456333482721,0.00208773865490808,0.0142309413418436,0.000951194240701225,-0.000124167412233311,0.0217161106790407,0.00310765801925594,0.000785900672522821,-0.00154803023238326
"122",-0.000132920054864427,0.00206897318427446,-0.00208338908298633,0.000228606353713801,-0.000238252434761166,-0.000619296028975924,-0.00390614505051312,0.00898523256849959,0.00926659366315663,-0.00310073611494466
"123",0.000332020330312766,0.00593609782977578,0.00974249412641681,0.00350682506350264,0.010320003979873,0.00520638854453614,-0.00128975629337424,-0.00230310842972414,0.000155539988934361,-0.00077756390523942
"124",0.00904066890841548,0.0116307767585364,0.0179184914926691,0.0202842756365429,0.00525754830938197,0.00152332023562596,0.0251870990603649,0.011080236238143,0.011669519760519,0.00622568534584866
"125",0.00362366936199909,0.00608673296331785,-0.00203103199143273,0.00796712386485821,-0.00609790864207471,-0.00296817888646328,-0.0046614344872814,0.000456887969964903,-0.0043063520904193,0.00116001076655725
"126",-0.00105038099032806,-0.00344534625923221,-0.00271367955502955,0.00443257108787187,-0.0112063371024914,-0.00557828478648292,0.0160755192610329,-0.00654184200317254,-0.00494284846904058,0.00926999570093279
"127",0.00525708979776263,0.00758872253194354,-0.00476193484436693,0.0171356774272342,-0.00405656613176686,-0.00236833105423684,-0.00211755918759216,0.0124041656952312,0.00838250569334065,0.00841948881502264
"128",0.000784165022412964,0.00343094048306103,0,0.00968938591894619,0.00359397290639185,0.00362445583820747,0.00374515479205262,-0.00862187604070552,0.00646548655273227,-0.0022770415146578
"129",-0.0142386321497765,-0.0146773520504691,0.00205069945502645,-0.0196936939905863,0.016949348940186,0.00684722925156267,-0.0304722940059292,-0.0122063099249407,0.00351795672306299,0.00722704709078603
"130",0.007089687530758,0.0131183953364196,-0.00341087289682829,0.00825485644868862,-0.0103274738065016,-0.00346271839339318,0,0.00447930672792429,-0.00259105315361896,0.00226594368689348
"131",0.0157904101652069,0.0167086055796781,0.00684486125007022,0.02195327267391,-0.00343966274384555,-0.00285350903075254,0.0125718173959442,0.00830393358407311,0.00886300400785434,0.0026375300692274
"132",0.00297928822441063,-0.00246510614418416,0.00475852942747013,0.01240696945607,0.00273657317314879,0.00224079171505354,0.00950176398610769,0.00732044809283461,0.000151499552476508,0.00150315505542631
"133",-0.000129295905350491,-0.00230627184353971,-0.00202982463050805,-0.0098040106308529,0.00961333529709352,0.00397241997798936,-0.00552157381456642,-0.0040880759013282,-0.0031803574614625,-0.017636035275769
"134",-0.000516102377158045,-0.00132115881073724,-0.00542376364150687,-0.00077765449998457,-0.00211691515636869,-0.00210286587079855,-0.00643609617000884,-0.00881734388375843,-0.00106350653296861,-0.00611145817995895
"135",-0.00180953318968713,-0.00727521036742329,-0.00477142124794239,-0.0122442676418265,0.00376995451107898,0.00359534108028847,-0.00546151791489446,-0.00153344991013771,0.0132319847908744,0.011529517868204
"136",0.00388415594610358,0.00441374469325995,0.00479429685783872,0.00995981270336532,-0.000233785953827392,-0.000123065092459185,0.00332025801721159,0.0015358049901617,0.00585408259438247,0.00341949609782533
"137",-0.0101245386130024,-0.00920308670405623,-0.00408998492604473,-0.00688185686013554,0.00903855041534829,0.00493970803602828,-0.0160382545515589,0.0007670632748773,0.00850619285162812,-0.000378725846339356
"138",0.00306188619168712,0.00317977001347347,0.00616030966219117,0.0289327704335633,-0.00162917979721944,-0.000368361446894894,-0.0174647877306542,-0.00766254063832905,-0.00162771525221317,-0.00454541746867632
"139",-0.0173412036940747,-0.0212710864938159,-0.00340136104392641,-0.0342291787135595,0.00372930836320062,0.0027055917150558,-0.0256747491853659,-0.0200774394506253,0,-0.00761027412690252
"140",0.00204906829414764,-0.00196058377504882,0.00068268240673941,0.00575122444209208,0.00197315637137763,0.00134861945233511,0.00135126899275173,0.00315237138009361,-0.00844818425302818,0.00881890096296867
"141",-0.0236789865621061,-0.0379161408564341,-0.0177352974068611,-0.0509650184618035,0.00834181198777117,0.00795923425455181,-0.0229421042632333,-0.0416342608348163,-0.0186846033278145,-0.0106421866674594
"142",-0.0196597574128496,-0.015178253230312,-0.0097225180956142,-0.0129546724358921,0.00287193392851126,0.00194482302488841,-0.0276239133178736,-0.0186885671431181,-0.00365571961444877,0.00960418518193684
"143",0.0156430158494285,0.0208199764207122,0.0168303388629123,0.0327355374577747,-0.00286370954391069,-0.00254654088541173,0.013494066735489,0.00818594005935203,0.00550363825080957,-0.0114154519572044
"144",-0.0112628260695751,0.00573942092451851,-0.00482744711235439,-0.0204668725553647,0.00723865627453701,0.00413309964687736,-0.0133144013155935,0.0122620161035778,0.000304150842518558,0.00808306373567436
"145",0.00487208839835551,-0.000527178612722223,-0.00762292742032877,-0.0039221921160435,-0.00216449863936019,-0.00277123880628505,0.0156249477590655,-0.00965819512601684,0.002127967743913,-0.00152730162096215
"146",0.00799012388336684,0.00368884645434897,-0.00488838477162845,0.0110561991536857,0.00252500219309182,0.000731140781434769,0.014685054448794,0.00495875866001194,-0.00060671924768696,0.0015296378393137
"147",-0.0257448827985178,-0.0175021880251754,-0.014034960247017,-0.0431427167911601,0.00663983969279913,0.00645491187525904,-0.0368021289686974,-0.014967222035067,0.0121414935823569,-0.0110728958450327
"148",0.016759100354935,0.0115795236828584,0.0149463388018027,0.0178470188011743,-0.00727827078534704,-0.00399349897920609,0.0260444582170491,0.00100202051480136,-0.00254918270957627,-0.0138994995789665
"149",0.0106694920080848,0.00255329064627996,-0.00210349757612605,0.00746004547333357,-0.000801767871318138,-0.000121661749748592,0.00404489041446232,0.0158463548225956,-0.000601232739081525,0.00548151681725861
"150",0.013941148551057,0.0209030167247053,0.00843281046873101,0.0335877834855018,-0.0121534071987132,-0.00692544475686807,0.0362550178746777,0.0279147526460752,0.00436212375020517,-0.00155763343848836
"151",-0.0296337416960801,-0.035185786533353,-0.0160279536862059,-0.0413587786930516,0.00139246815923744,0.00562856292572844,-0.00174285966108279,-0.019009535488116,-0.0196195605640062,-0.00780031722738583
"152",-0.00467724001702996,-0.0141775569364661,-0.0141642867607384,-0.0173345508096689,-0.00231742591479722,-0.00146076328714917,-0.0331676260909671,-0.00749061640206938,0.0169569357921926,0.00353769611988386
"153",0.00359303737643502,-0.000181205967607068,0.00143665773391533,0.00987861424455505,0.00290346324259461,0.00158409459624531,-0.00416677116325581,-0.0045942888291598,-0.00465672224725844,-0.00705053381947773
"154",-0.0152859445068955,-0.00986045378495271,-0.00286934834296548,-0.0258519273506386,0.00266423115224534,0.00364938643641155,-0.0376566300568827,-0.0214275718173007,0.000452746741540944,0.0031557362828909
"155",-0.0137751178411848,-0.0244859259914867,-0.0165467570170523,-0.0392896385546739,-0.00358085756300386,0.0018185514339959,-0.010869661568372,-0.0296443649644578,-0.00241369735384378,0.00747162273480795
"156",0.00751566405203508,-0.00290334529023584,0.00219453294619432,-0.0170048335887028,0.0103183167847538,0.00387095476227417,0.0257873194047358,-0.0218713888430772,-0.0219264640220684,-0.0171741360556121
"157",0.0183673362161205,0.0186920899897556,-0.00729915928254421,0.0316452335719222,-0.00401560492069775,0.000723865261023082,0.0262823672722414,0.0216510562969028,0.00510207173778587,-0.000794281750049253
"158",-0.000483876719418741,-0.00138289062661601,-0.0110294813218508,0.00204521102440292,0.000575904189412224,0.0021674843145203,0.0167013020309696,0.00052109566633729,0.00169206270751987,0.00278215339106791
"159",0.00200506806658307,-0.00277031012664364,0.01263941698912,-0.00367350978253256,0.00483644840158681,0.0043276973291857,0.0150584848858806,0.0111106507866325,-0.000767859301235019,-0.0015852880109033
"160",0.0118677984304822,0.0247223731783011,0.0132161470204983,0.0430151232475411,-0.00160436132662678,-0.00323132897325484,0.0080914422691849,0.0317652141376399,0.00507149223912728,0.00238181403621773
"161",-0.000886235107046107,-0.000813248730227367,0.00724608552873685,0.00510597711112393,0.00344340237887586,0.000359836339017816,-0.00709036749647762,0.00931925099859354,-0.00137620790898463,0.00316823425738266
"162",0.012353015805183,0.0215227090678038,0.00503591452020791,0.0238374402546291,0.0049186089509563,0.00035995509123854,-0.00633247030463124,0.0189612733440492,0.0122493190093194,0.0118436731577627
"163",-0.0093035788897764,-0.00894096263319188,-0.00787384550626125,0.0045799816059402,0.00523655551454283,0.00275969920534025,-0.0135591711233048,-0.00728159206840728,-0.0019663893213373,0.00117050424605614
"164",-0.0219805198351637,-0.0241179937537898,-0.00937954578849232,-0.0406533455393291,0.0016987549859695,0.00514349279865978,-0.0316152665979671,-0.0221675900915345,-0.00591098790947309,-0.0105221384053501
"165",0.0196216625536725,0.0259040417955128,0.00946835465451601,0.0396038748393359,-0.00271328689173889,-0.00380903485469464,0.0262596090476932,0.0218371201124339,0.00731825017949372,0.00945246275909684
"166",-0.00266119555574829,-0.00562117799519191,-0.00649363614931553,-0.0051041657063744,0.00668763713510456,0.00501866219513492,0.0048409669510503,-0.00897267861170081,-0.00408652943847421,0.00195096581230558
"167",0.00985285195521013,0.0171376710395605,0.0217866090869918,0.025807399489532,0.000788163430373245,0.000237842036632019,0.019958733468574,0.0139921373222889,0.0109421575558286,0.000389366640277888
"168",0.0100951600133397,0.0096154526604344,-0.0056858043796042,0.0168718368267584,0.000473704586966495,-0.00186123549835882,0.0134951276810902,0.0159091950072008,0.0138305027283752,0.0112884887874316
"169",-0.00865291605204421,-0.0139799052979107,-0.0192995755588122,-0.015123654048729,0.00801776916372599,0.00621542451152068,-0.0239680972592975,-0.0209334067012434,0.0017793000658568,0.00192459985923144
"170",0.00230084836120947,0.0022154627599511,0.000728867562922009,0.00782722602579722,-0.00257638075210398,-0.00213786439435315,0.0061394497706857,-0.00522274897555408,0.01924220009598,-0.00384172346283407
"171",-0.0139066499090779,-0.011582737103802,-0.00509842432501229,-0.022559496210091,0.0141513503737123,0.0107153462304257,-0.0187121262631141,-0.0164069147534379,0.00769674691117128,0.00655603403984628
"172",-0.00191686389495593,-0.00581456687079573,-0.00878478403871175,0.000756857898968732,0.00775246783574279,0.00223734014761057,-0.0189300428131013,-0.0145120105037594,0.00331465633830019,0.00689651548866221
"173",0.0116600427682814,0.0197051411459188,0.0103401193262109,0.0201885812228639,-0.00077001034085511,-0.00211504745031821,0.0180278941896934,0.018957062850707,0.0129272329965284,0.00228314746503155
"174",0.00257696233544058,0.00326465691225564,-0.00292446782040079,0.00355822685076679,-0.00373947990504198,-0.00247323832903612,0.00179861091369005,0.0101329952503719,-0.000850794137158162,0.0106301868737808
"175",0.00703304992491693,0.00562862961704402,-0.00733126772577464,0.0110782830095528,-0.00894098134072308,-0.00590428444240931,0.0183679024433021,0.00970233910337681,-0.00539308835357777,-0.0075131534517725
"176",-0.000067195786397134,-0.00997017842272074,0.00295436537915239,0.00197196311811743,0.00144768277599083,0.0013070349105293,0.00474587118317027,-0.00716644733417116,-0.00128430361631549,0.000757043374380428
"177",-0.00537276097706851,-0.0167841639439079,-0.00515476225446776,-0.00634228566320272,0.00478282845793876,0.000592161315494,-0.00188940026231954,-0.0247700015832637,0.0140020435491368,0.0117245866427997
"178",0.0294396847835368,0.0420485480912887,0.0103629201800133,0.0484228587790974,-0.00752701166471281,-0.00106574798951187,0.0311022476771026,0.027754310310224,0.0102859798466115,0.00373824050057459
"179",0.00590301997141274,0.00353475590999852,0.0109890785472468,0.00454826576858802,-0.00925774259672496,-0.00356027647740176,0.0203275638184566,0.0193127761469973,-0.00376564869312324,0.0085661949880711
"180",-0.00704199962566199,0.00223388420100679,-0.00362327750789471,-0.00313463830739302,-0.0189120155838297,-0.0113146633066039,-0.0122105745921655,-0.00851018409565873,0.0180596528069437,0.0155096524025742
"181",0.00269863161491624,0.00642961574587742,0.00218160726626504,0.0132773672502382,0.00849045134281079,0.00505863151356678,0.000260204549973553,0.0131568700741951,-0.00522559123727184,0.00690905679580123
"182",-0.00184255885193474,-0.00170336481528877,0.00362869406709243,0.0124140146200282,0.00284516780734667,0.00131869417590269,0.00858579039441687,-0.00145187249113188,-0.000829375218654893,-0.00180574604944927
"183",-0.00197766324380866,-0.00392520643456329,0.00578422725780925,-0.00374653918449008,-0.00351697241493842,0.000120265888877036,-0.0165532814946034,0.00226160943029763,0.000691795803704931,-0.0072358181019565
"184",0.00528447587401115,0.00436879999066475,0.00862698698024911,0.0133330635247786,0.000910527632447922,0.000359094166186846,0.00569019207600774,0.0169250447707769,-0.00456244975632647,0.00145768792851686
"185",0.00591342781701143,0.0119403047501434,0.0228083244847279,0.0148449382338249,0.00693928522684395,0.00323003013980605,0.00947352923390299,0.0112536391858253,0.0097221805555554,0.0262008927706412
"186",-0.00333146622497538,0.00463533091222179,-0.000696868486341984,-0.00631664442333868,0.00225955224308683,0.000357547480760889,-0.0032589093476173,0.00705288403263893,0.011141747364859,-0.00319145367419116
"187",0.0112725034799659,0.0100671280703544,0.0111574345497361,0.031448650768783,0.00571409021321201,0.00119657254314776,0.0265466962329173,0.00498086652666285,0.00530540048142014,-0.0103167347210077
"188",-0.00136028994332638,-0.00298998201771672,-0.00275853208823684,0.00681171814300674,0.00314978419763534,0.00215117795103281,0.00917206430286743,-0.00263262852442792,-0.020974343140072,-0.0201293040553866
"189",-0.00201227272373161,-0.00366544633910704,0.000691588665405085,-0.0302839143490033,-0.00291605505367232,-0.000715340614004689,-0.000252544554585676,0.00155242407057021,-0.00621970991623244,0.00110047505025279
"190",0.00156125053170331,0.0052676389083961,-0.000691110701077635,0.00996709407336138,0.0038247300683083,0.00178968888322517,0.000378987775617956,-0.00465110074952335,0.0134909731991384,0.013924485602435
"191",0.0118812803020723,0.00756862517602341,0.0131397365843875,0.0333551385126516,-0.0107575095894195,-0.00881579930084275,0.0198156556639584,0.00934579294627991,0.0072732122708985,0.0028913363212475
"192",-0.00532591670424531,-0.0114741447156635,-0.00546078535327499,-0.0106320653164975,-0.000793407983270655,0.00360579812799444,-0.0111384421342122,-0.00925925783967396,-0.0118529015843896,-0.0209009532259744
"193",0.0094182257913884,0.0125260359748325,-0.00274551168299308,0.0155726125918589,-0.00124641992661079,-0.00311347506469573,0.00575702196092975,0.0171339537348463,0.00772090180230101,0.00699301195640767
"194",-0.0016613466833586,0.000412400805846813,-0.00206464345225976,0.00133064817366657,0.000567215586389835,0.000961664568288612,-0.00136915274061822,-0.00137779149213157,0.00369414440794325,0.0116958755188288
"195",-0.00480132176572989,0.00412203349426421,0.00137948945528032,-0.00879546987914048,-0.00102066196511319,0.000119825737218582,-0.00672874725430128,-0.003987335471755,0.00749731451066915,0.0111994302013048
"196",0.00553205881039642,0.00615775511616712,0,0.0182580415231384,-0.00488344023893839,-0.00335995640619313,-0.00727625012288979,0.000769761450125195,0.00920027010146018,0.00464463410506832
"197",-0.00844406342829129,-0.00873138143511731,-0.0117079986242382,-0.0122254371698546,0.000228340476359223,0.000962727342953995,-0.0205991934302905,-0.00846171902843795,0.00737368319472775,0.0170696735864164
"198",-0.00793492021141096,-0.0113598956092915,-0.01811834414863,-0.0185340377890293,0.000342601952121102,0.00276688453804486,-0.0166454863573657,-0.0217223544621982,-0.000266116585921239,0.00104887679717081
"199",0.00305657294169448,0.0122397442436084,0.00141930187488248,0.0230872519793472,0.0109485324938143,0.00611837551851457,-0.00275507743053927,0.00475847482491232,-0.00825350073535003,-0.00523930066369616
"200",-0.00363019703637868,-0.000493289544029607,0.00425239570472646,0.00505723734342167,0.00552764844519782,0.00381521683380659,0.00263148112884104,-0.00552476553110881,0.0201342281879195,0.0179073168434274
"201",-0.0261569452529566,-0.0198337982160064,-0.0197599831182678,-0.0427675236344222,0.0149225165490419,0.0085521154213315,-0.0322832263878455,-0.027301964609576,-0.00394740789473691,-0.00275953735000611
"202",0.00581297431307082,-0.00503794215435471,0.0057592413702281,0.00722730678607397,0.000110335783753079,-0.00188434054993547,0.0123404071071422,-0.000489445835774038,-0.0145310309589576,-0.00276717346854638
"203",0.00810411413630918,0.0156118149927293,0.00286325268596954,0.0277237026581909,-0.00132585310469446,-0.000235624005499591,0.00870732579360545,0.0179588551928092,0.00844510746501625,-0.00693725997684724
"204",-0.00184543670719639,-0.00124632878962905,-0.00428248468630033,-0.006537557750949,0.00741582791480422,0.00507457848444282,-0.00398442475782002,-0.000160040765461389,0.00385476523243011,0.00349284216203993
"205",0.00237690200869478,0.00582381994565973,-0.00358431825157945,0.0127138565139182,-0.00340633007524094,-0.000821830221945263,-0.00266656870456372,0.0131539059942438,0.0067532047174208,0.0233204754837524
"206",0.0117226756146891,0.0168732486453387,0.0172662304517246,0.0283261476465728,-0.00231508566173844,-0.00246790445871603,0.0147060122481957,0.0186825632220284,0.0218335265268121,0.0153063169226604
"207",0.00332029700567649,0.00618191373908705,0.0134369248248571,0.0230063620750971,0.00386721621245623,0.000824718384696332,-0.00724652963117578,0.00326394644570782,0.00553483059506155,0.0164152409450689
"208",-0.00694252745531132,-0.00727584797547476,-0.00488488849428359,-0.0188906446994888,-0.000550651125708623,0.00105904357158848,0.00451249639941764,-0.00325332775813503,-0.00985669444994774,-0.0224126033472398
"209",0.0103879222746945,0.0146581506485803,0.0070126898724332,0.0219438828213059,-0.00902993293800747,-0.00670278660609458,0.0179676636363413,0.0219147336994612,0.016418940308182,0.0283210275855652
"210",-0.0234074687764573,-0.0244780762671079,-0.0125346631326069,-0.0403734363716898,0.0129931473825211,0.00816192856801656,-0.0356907898662565,-0.026768181289057,-0.00877643059871147,-0.0127869289061899
"211",0.00112552260543941,0.00822700961820999,-0.00282093566189301,0.0056720710493332,0.00319511210899104,0.00270971891871774,-0.0197846248869123,-0.0078137199719136,0.0243808802771717,0.0215875633978628
"212",-0.00760529803932841,-0.0134639201049574,-0.0169731678245698,-0.0347694012137114,-0.000439372063361976,-0.00117467132324323,-0.0142795019741565,-0.0195305948681092,-0.00100215455337194,-0.00650202454672566
"213",0.0134617011004372,0.0140611657329115,0.011511042258094,0.0379479737033666,-0.00483555835795835,-0.00176487327558261,0.0104467411791918,0.00883533995538044,0.0210658307210032,0.0261779946862162
"214",-0.0273559129716343,-0.0160684799260115,-0.018492135996615,-0.0318587949632806,0.00176722876205049,0.00365381478888627,-0.0337747286934746,-0.019586256263014,0.00994716934790607,-0.00510201048791581
"215",-0.00507061410097376,0.00886997780215637,-0.0159421929981683,0.00511176510803568,-0.00176411117404429,0.00223089582889502,0.00627791307907133,-0.0035727948149521,-0.000121534536029588,-0.00256400139839019
"216",-0.0137262806312005,-0.0230073339780787,-0.0132549828554372,-0.0235219789804773,0.00850244350290841,0.00597680292973846,-0.00340298570595832,-0.0203749252337623,-0.000608087050659512,-0.0003214058130524
"217",-0.00992148730081543,-0.015979817797096,0.000746457658829192,-0.0553385870666256,0.00361285043922388,0.00174652640967277,0.000142690098884346,-0.0257904095710222,-0.047213397420297,-0.0218579729895122
"218",0.0304798617043007,0.028632311515161,0.0171511187903453,0.0706407895591592,-0.00370838836396215,-0.0051151727554869,0.035846511290033,0.0401366964163938,0.0104725411057773,-0.0190600112852922
"219",-0.00276861966598441,-0.00290804181772786,0.00293304541733952,0.00096558964554494,0.00109462511834035,0.000701000482944636,-0.0146938608480721,-0.010673199746856,0.0146612229021277,0.0224454312693505
"220",-0.0144241668674087,-0.0166667297337182,-0.00877209540838042,-0.0230221190722709,0.00940741601746531,0.00560640029717874,-0.00557515612480541,-0.0182571906366428,-0.0290234433112039,-0.00982962716745794
"221",0.00171793536551945,0.00423720823736984,-0.00737497268596066,0.0123746246203704,0.00140865129929635,0,-0.0190607484807915,-0.00422667563616963,-0.00256570888642882,0.00330906930670882
"222",-0.0139242669338624,-0.0270040189205014,-0.0170874120479615,-0.0460986859943814,0.0064930679537285,0.0072003050229501,-0.0191456360340448,-0.0280135766728004,-0.00655951125401932,0.00758579294261863
"223",0.00612143075086236,0.02228948965563,0.0264550524892304,0.0274693946399389,-0.00107508539123635,-0.00265219778169024,-0.0233065052267406,0.0155462578315058,0.0288710908563203,0.0248772327886559
"224",-0.0204645233500647,-0.018494799601682,-0.0176729999848465,-0.0503519761954589,0.00581167736896382,0.00786221937129494,-0.0074573131323844,-0.0223603201521001,-0.00138417010967451,0.00127765068033292
"225",0.0172923831257001,0.0215228188000596,0.0224884324621055,0.0295495738870151,0.00299668371727391,-0.00298246256953549,0.019083469244362,0.0362421913556661,0.0238155112926473,0.00925023354463761
"226",-0.0220632795565719,-0.0197158845569588,0,-0.0396933746377771,0.0197374012684308,0.0136916717327058,-0.0375999312439347,-0.0290325288115001,0.000615421538461502,-0.0123260774232595
"227",0.0114930166689913,0.0125164099605324,0.0161292956574379,0.0382955373682154,-0.0095218752918349,-0.00930664178507157,0.00735416774610154,0.0307747592198213,-0.014760208557434,-0.00800003976861519
"228",0.0319848035949026,0.0323956301100772,0.00937954578849221,0.0547810760086909,-0.00675970336012954,-0.0035526042996411,0.0468443008510928,0.0154369513809964,-0.00661670428506134,-0.0122580734124823
"229",0.000339587059499102,-0.00908330616085762,0.00357413595901068,-0.0122585678971143,0.00861480204797527,0.00563453922694035,0.00799077051335062,0.00133637178115231,-0.016212152821415,0.00228622915887211
"230",0.0100557161485935,0.00374999211661864,0.00213654535236074,0.00849148070288686,-0.00485071629311762,0.00137155981408776,0.00922415900676321,0.0060063102224257,-0.0122636562629492,-0.0123820652419223
"231",-0.00659292093207786,-0.00356983076805573,0.00142158265998504,-0.00867874392603918,0.00793599631038355,0.0039529320850118,-0.00728295594533102,0.00364817255104222,0.0124159208484222,0.00725844226775885
"232",-0.00893791619327611,-0.00599909788798181,-0.0106461544821596,-0.00261355893755921,-0.000105409134551704,0.000913179828276212,-0.026183780631134,-0.0133840751440543,0.0143076522011707,0.00458558632946859
"233",0.016739719748591,0.00813040333435544,0.0186515056515189,0.0444126033917824,-0.0119275346011029,-0.0037624018134339,0.0285125778198929,0.0217719617400531,-0.00969779572549634,-0.00749915544072055
"234",0.0143133961906641,0.0106432427448735,0.0126760713019587,0.015742584207568,-0.00875958825503553,-0.0052645576153092,0.0359094411057561,0.0136044095319876,0.00941124288736761,0.0180682734706157
"235",-0.000198597122705868,-0.00255070820462977,-0.00904036936596753,-0.0118555680411088,-0.0112075208482618,-0.00644253470804135,-0.00485318975269022,0.00258700659191069,-0.00970146114269388,-0.00322681525340973
"236",0.00775276636141209,0.0112176139197737,0.00280707865154928,0.000312549587313304,-0.00599524800515405,-0.00231616781903643,0.0250802522374853,0.00403248265779599,0.0178117307331229,-0.000647459196076228
"237",-0.0274195474123864,-0.0268355498942128,-0.0216936066555369,-0.042354014034613,0.0196278789972872,0.0136948518351891,-0.05722449085212,-0.0224903073603734,-0.01450005,0.00874629264896143
"238",0.00987121437271021,0.0233846666609323,0.00786863237999857,0.0300066149543305,-0.0103241610399734,-0.00835722837930397,0.00317164805695458,0,0.0209284891389392,0.0272961382131933
"239",-0.00207544709820473,-0.0197377635220541,-0.0205819026015447,-0.0274857091115677,-0.01086643946495,-0.0073898876894023,-0.0172466021903745,-0.0164331059277806,-0.0247235439116299,-0.0106282956909713
"240",-0.0126797006158279,-0.0252318601554168,-0.0391306727338105,-0.0238343775971503,-0.00461389589897576,-0.00290774037934782,-0.0302714584562116,-0.0342525768703734,0.000254738853503245,-0.00695106564738879
"241",-0.014269284274001,-0.0173995901903597,-0.0173454164028385,-0.0426284259585809,0.00893925535617202,0.00594955291960919,-0.0180972982567528,-0.0501731684652021,-0.0049668876069876,-0.00489079563714301
"242",0.00558376072456768,0.0109909897206337,0.0176515905918262,0.027454268985033,0.00645410017976911,0.00197107683789643,0.0129011769162997,0.00273195060093023,0.0143351215026926,-0.00425944207669848
"243",0,-0.0101811177686408,-0.00678728020324915,0.00651106483369035,0.0132600325455601,0.00798536606509126,0.00833993208083994,0.00999153274618991,-0.000126208201892797,0.00954259968372395
"244",0.00630683447866875,0.00392258544060597,0.00379657790040611,0.00545772135762856,-0.00214512749555318,-0.00160588062015321,0.003759444896001,-0.0062952114866569,-0.00719333688019519,-0.00423733058600284
"245",0.0144151038876232,0.0145869754182106,0.0151285469309952,0.030156914823759,-0.0146193425122731,-0.00724604852020183,0.0170786331113826,0.0130323695503434,0.0181771963436428,0.0117839818799261
"246",0.00742604009541181,0.00679760192471512,-0.00165626104792826,0.0169130397227275,-0.00469100172574921,-0.0028966109494476,0.0272501883800946,0.0189192180827122,0.000499388277138246,0.00744093606279606
"247",0.00214427969945241,0.00550262562504544,0.00452501535372996,0.0051835119193544,-0.00876749970842361,-0.00476292545005663,-0.0166330137132936,0.0150307645577412,0.0172198404943829,0.011881835103565
"248",-0.0125712427840621,-0.00277978675360968,-0.0157660165355747,-0.0230758601665397,0.0109008147380112,0.00671309096758166,-0.0194550659697155,-0.0243899860432898,0.000490689419431423,0.0034910490379898
"249",-0.00250577822072418,0.0083624525487922,0.0114417759386638,0.00376094765739921,0.0155946993752787,0.00803104715934544,-0.0147412984944172,0.0157143024013324,0.0176557385398661,-0.00316255885803629
"250",-0.00739961609475115,-0.0122668878140141,0.00226242707985747,-0.0120291410627522,0.00605528297785884,0.00461837627992989,0.00305355585215517,0.00123034978734649,-0.00650603614457834,0.00126896397825904
"251",-0.00875454142622212,-0.00271119821872268,-0.00451489284875173,-0.0165006213425194,0.0144022975723586,0.00712587650716134,-0.00837154213759228,-0.0043898632550694,0.0291050452231998,0.0275666024282257
"252",-0.000483053708982717,0.00175388701728818,0.00377924767754068,0.00899762963804607,-0.0013770533259424,0.00205461267017837,-0.0323867391894161,-0.00370356753840073,0.00836670977649412,0.00770883958221713
"253",-0.0245066269187432,-0.0234611084142807,-0.0256024539278635,-0.030036753377831,0.000211103814771185,0.00261901321136349,-0.0317256465965057,-0.0219506570349396,-0.00514202407385755,-0.00581387407030654
"254",-0.000848823548182609,0.00502019914042906,-0.00618222739996965,0.00732694392373512,0.00434965671713239,0.00181627048721067,0.00933804641446678,-0.0162897587377726,-0.00422882664967084,-0.0181595601336975
"255",-0.0161482734553615,-0.00909849370325122,-0.00233260850879746,-0.00775389796048764,-0.00116172418272886,0.00215504743219563,-0.0363577497497656,-0.0220791884382113,0.0237112430238733,0.00909093024415042
"256",0.0105099906164954,0.0041410483757276,0.0218236838284818,0.0327800400857994,0.00190358786180478,-0.0015842441169589,0.0197069713460403,0.00564459743542045,-0.00265033420892291,-0.00994093566611409
"257",0.00655402068506583,0.00080677716055777,-0.00839053631259068,0.0117850219463849,-0.0135094005727793,-0.00271983428695,0.013214367248604,0.00187104532115012,0.0196417901915036,-0.00470664262171938
"258",-0.0080683877485207,-0.017377589944241,-0.0169230427386049,-0.0281269593222061,0.00781040091444485,0.00636337254668518,-0.00163025314234433,-0.0252099891132497,0.0037393994334276,0.00914241888765055
"259",0.00806276515993543,0.0165908968899482,0.0125193210571037,0.014708622955947,0.00371542211825671,0.000452027075156236,-0.00277624723856951,0.0153253247211822,0.0108376493376012,0.0124962089895626
"260",-0.0220129641316857,-0.0312949109852088,-0.027820566035198,-0.0452318405067965,0.0112115189217041,0.0065455030151671,-0.0260352251805488,-0.030943294128266,-0.0173107324401304,-0.0123419810154484
"261",-0.00861251334190094,-0.0216603720916457,-0.0182827708821331,-0.041610809318769,-0.00721719719511593,-0.00190657582636777,0.012945110768404,0.00272555127984253,-0.0146607686023587,-0.00937191995711351
"262",-0.0259166183443298,-0.0142873891425744,-0.0137654116735858,-0.0291162017005472,0.0129575590373636,0.0080877997865807,-0.0121159676941429,-0.0108736043301751,-0.002306770552714,-0.0129297788189532
"263",-0.0102674264923376,0.0010560883410855,0.0262725516921734,0.0228132783682657,-0.00686361108145328,-0.00144703855775352,-0.00840079751857703,0.00706708724023963,0.0106358150289019,0.00383388391305206
"264",-0.0101465694560247,-0.031258942464217,-0.0367999289834803,-0.0251112450738022,0.0106817390972032,0.011158511149197,0.0337174774959583,-0.0183234736199698,0.00857927267397107,-0.00350091581404965
"265",0.0240208032286362,-0.00653284015322619,0.00332222711888552,0.00636356695531459,-0.00227948159263824,-0.00463513688631922,0.0817903288277588,0.0127084896413487,-0.00317567206931324,-0.0188438187034397
"266",0.0084416966815708,0.0297897043501394,0.0165561829167438,0.0194219978986223,-0.0200446140972894,-0.00909160915297447,-0.0195460644910043,0.0284313842903927,0.0249175449416035,0.0247395512072714
"267",-0.0144457221095226,-0.0201239952895084,0.0154724206090635,-0.0152118427739741,0.0168508058294035,0.00928702000445081,-0.0139076786997623,0.028599197606576,0.00244228458165452,0.0222363674138357
"268",0.0165367523522588,0.0156992217248368,-0.00561322864604885,0.0247449009786604,-0.00375157838700724,-0.00365914448484506,0.0371414484908741,-0.00185428823784717,0.0160575520689628,0.00466139951663203
"269",0.004953696140793,0.00767943970991158,0.0169352862768217,-0.00490255606973733,-0.00679996705899377,-0.00400519286574341,-0.00604443564879276,0.00185773301031733,-0.00653948773841961,0.0083512203980638
"270",-0.00735747263565423,-0.00347276714285338,-0.00475816727830214,-0.0131626911238178,-0.00653027620705693,-0.000446584117021032,-0.0234112406241844,-0.0157562276004234,0.00998349950667032,-0.00858889055647272
"271",0.018234125636295,0.00948685953623674,0.0135456560549425,0.0200448489481926,0.00710294046364734,0.0051412047251751,0.0238170148353984,0.0169496676109782,-0.00716919415966089,0.0049505395663092
"272",0.0160879673114189,0.0138090430653977,0.00864815504745353,0.0199428319599664,0.00601167768947075,0.00324503693901113,0.0389235124230327,0.0203704115191787,-0.0224289272991482,-0.0175493094837592
"273",-0.0126091195721454,-0.00813447130325506,-0.00311818590736745,0.00307993535746265,-0.0102918003932478,-0.00555904098124826,-0.0155130279145859,-0.00381146851172398,-0.00279798551310539,0.0175493516543039
"274",-0.0267740387328466,-0.0500670082112697,-0.0336197322485399,-0.0538380421675838,0.00763959679817039,0.00704414153554911,-0.0316634472252899,-0.0435418933961362,-0.0159371271815292,-0.00831537447744168
"275",-0.00805217756322607,0.00552154921732795,-0.0129449088258343,-0.0163762741774102,-0.00305300482662385,-0.00177629168673932,-0.0191895425106859,0,0.0144844548357663,-0.00465840677163776
"276",0.00661402812129386,-0.0108825995384734,0.0057375304571663,0.0169561641308029,-0.0215468152359146,-0.0112334647852058,0.0241041889876048,-0.00857127577429617,0.0101180554283773,0.0121684457745848
"277",-0.00642100233915111,-0.00353279500493153,-0.0252647639919378,-0.00188668295032812,0.0114424728563221,0.00843628732127133,-0.0310256273233656,0.00192148525309954,0.0127991321713774,0.0299014221653737
"278",0.00510996101083849,0.000911867700279734,0.0100334248354799,0.0123962656630496,0.00416206201237945,0.00223165134054826,-0.0200315079519064,0,0.00362639560439559,0.00658490632753428
"279",0.00927124031545934,0.0254021170011045,0.0149005823190511,0.0161266890117528,-0.00595209078327263,-0.00211494249282385,0.0315464758937321,0.0134230903585739,-0.0218986089587516,-0.0202200517606466
"280",0.0102228185725128,0.0141135157712808,-0.00734077038202052,0.0224833943454437,-0.0105835630345888,-0.00423848864639054,0.00468095853426909,0.00851458115311976,0.00123138920337218,0.00819414455935585
"281",-0.00879963928466954,-0.00778586590759889,0.00986029183296444,-0.0128626549410353,-0.0146974229407947,-0.00548849552684771,-0.00745435643971537,-0.00093815527673069,0.00301874993249651,0.0201685945015921
"282",-0.000222062153156788,-0.00392297494988181,0.0122047091697532,0.00713417995751264,0.00767629860987706,0.00214052719170854,-0.004068336355457,-0.00187825747967396,-0.00624230304583995,-0.00472116848927839
"283",0.00281200363149603,0.0125058790477528,0.00964655567852368,0.0130825708005551,-0.0101217312198769,-0.00719292818253414,-0.0174392812848401,0.0169329767629849,0.0272574306840732,0.0326120194826895
"284",0.00295155629131361,-0.000486405181475913,-0.0207007420456533,0.00834783968555097,0.00692765661271477,-0.00090542390858106,0.0233451586040103,-0.0129507650824301,0.0181261843606424,0.00516786232688937
"285",-0.00831368924532849,-0.00136200102006756,0.0073172705598239,-0.014010018051427,0.010592296075784,0.0103101915777664,-0.0226561664855565,-0.00674802827200005,0.000107271559572464,-0.00542700647917216
"286",0.00615792586559527,0.00964636012342934,0.008070909832669,0.0134195033582138,-0.00572682816445269,-0.00280335352635597,0.0235013691445334,0.00490706858220835,0.0015013297587132,0.0137852753837973
"287",0.0126087841446771,0.0147653986846146,0.0208167839956797,0.0186231767989322,-0.0102151591635965,-0.00663604860398892,0.0309280489399928,0.0140844335623445,-0.0069600707459051,0.0096317030604518
"288",0.00750025753692785,0.0194958583947362,0.0109802736148663,0.0132081727129212,0.00032924602964135,0.0024909059967142,-0.000606293458736529,0.013888890409165,0.0104593597252396,0.0213242670851113
"289",-0.00101213346601559,-0.00335849936022303,-0.0054306860053781,0.00843919321173137,0.000878320761336759,0.00237228155559466,-0.00712552633352737,0.0100457903383904,0.0114182052226892,-0.00137369983327418
"290",-0.0097667568998262,-0.00393117729172265,-0.0109202262449559,-0.0107496794198139,0.0177647611745007,0.0117166810759244,-0.020766801044571,-0.00542546061920868,0.0127663959988014,0.0096287237141659
"291",-0.0222840445086936,-0.0247131833745603,-0.0118296889854613,-0.0397524866417223,0.0153005029874107,0.0106900766885467,-0.0174642876521308,-0.0334541138039408,0.00197939372808409,-0.0163487644500253
"292",-0.00239127221296842,0,-0.000797997699828801,0.00544371497876983,-0.00257804208469625,-0.00254220890592749,0.00539611986352306,0.00169300826023022,0.0110209814930338,0.0146813734667879
"293",-0.00382027777507077,-0.0112724045743262,-0.0231631224077775,-0.0232228729056457,-0.00971783601114018,-0.00376694804605848,-0.0080506174717706,-0.0159628390441048,-0.0211846775233376,-0.0035489822077398
"294",0.00631598628695063,0.0109137969914506,0.00572358203432644,0.0210032856277169,-0.0119706027734906,-0.00433776502033689,-0.000954797858569556,0.0160308482455345,0.0266862891363731,0.0219177486587276
"295",-0.0206976046030952,-0.0113749021461423,-0.00894291141741854,-0.0342856130867751,0.00534909380979709,0.00804276299597984,-0.0458747680744525,-0.015965394754294,-0.0124846601260268,0.00750686883795959
"296",-0.0103009345948708,-0.00887251452265436,-0.0147660213655113,-0.0138316512940448,0.00130236400529293,0.00343542926450158,0.010017091280659,-0.0112622497391703,-0.00424874611398962,-0.0101118449885799
"297",-0.0131832048626963,-0.0102314228956153,-0.00416342960610139,-0.0175500623634089,0.0147453115916776,0.00717791136476054,-0.0161984787655448,-0.0173743233014056,-0.00228944748837334,0.0188172265118327
"298",0.0359378976621147,0.0318061256580378,0.0292641685355162,0.0672567844552945,-0.00854829698324489,-0.0108555869334631,0.0710681958256392,0.0451867719598,0.00125164281052537,0.0155672258795234
"299",-0.00935148745872783,0.00250435735362586,0,-0.0185261444986151,0.0192910451602795,0.0115296856058777,-0.0214899754325888,-0.0203007926185373,0.0106261487785426,0.0109120036113952
"300",0.00220776932947375,0.00490080319363817,0.00324963246048671,-0.00911003574646352,-0.00782354324036172,-0.00526041204128103,0.0125040126093423,-0.00230195961050184,0.0137098646797265,0.00102792855388745
"301",-0.0154959246861192,-0.0253393735010571,-0.0663971103395585,-0.0354517705791066,0.0123611592256176,0.0103553654424231,-0.0163077041500862,-0.00576950328543779,0.00376248744203722,-0.00128365835410771
"302",-0.0101071511407212,-0.0171691275483581,0.028621161908867,-0.0247065751099471,0.00768368735564162,0.00501621317548229,-0.00676001718176789,-0.0348163773177921,0.00466010540634287,-0.0401027999348437
"303",0.0415430396107677,0.0303457622206078,0.0286678627915298,0.0519936385744126,-0.00386448419968644,-0.00683513765743249,0.0510453725793825,0.0320640107524293,-0.0269234451330734,0.0222280619906789
"304",-0.024769550002015,-0.0382677988427911,-0.0303279943231386,-0.0600519843822698,0.0165687128253944,0.00863028529720689,-0.0109469031656981,-0.0194172298379762,-0.0358549119170984,-0.0432275970356528
"305",0.0185226830478327,0.0126925981404644,0.0185967778783185,0.0168423545934808,0.00247540124469503,0.00216584296834088,0.041777064548308,0.00406240140074687,-0.0336414119342067,-0.0402519045767038
"306",0.0199877057692341,0.0179052478800101,0.0307053987962413,0.0383357446191968,-0.0193454343767854,-0.0176159266553061,0.017058218379252,0.0392700655161671,0.00211315750803442,0.0182596148216252
"307",0.000965156655560406,0.0177856852266034,0.0104670547039547,0.0153523204377171,0.0041975182734213,0.00352037146765416,0.00788435701770229,0.00954207934766793,0.0291898452650354,0.0100869355330777
"308",-0.0122357863406337,0.00384044669331907,-0.0079682090116997,-0.00811343356798022,-0.00417997276137305,0.000767346149161963,-0.0264204428659855,-0.00378080732059993,0.0115388759342541,0.0299583839720059
"309",-0.00315327284846778,0.00124356944104798,-0.00321291887650232,-0.00483313679604191,-0.00703062802812748,-0.00131401871098269,-0.00424482521290126,0,-0.00362477600347211,0.011042175200366
"310",-0.00956464598732643,-0.00487215870833457,0.00402906299077688,-0.00179383056447768,0.0097223759644034,0.00394814310048575,-0.0153777682716685,-0.0153700382196028,-0.0169056496565979,-0.0237079151963853
"311",0.0034977531163678,0.00806359197243833,-0.0072228430194281,0.00591402668351759,0.00355839272548231,0.00174796024878043,0.0066489307612323,0.018500847658026,-0.0159990536351454,-0.0240109860613007
"312",0.0351594080233859,0.0318067106490119,0.0291025061477415,0.0383985066607782,-0.0162747259084053,-0.00874311363785008,0.0491553161081912,0.0454119779377657,-0.0392655994130915,-0.00559131338682139
"313",0.000659126575671687,0.000368943089121387,-0.00157089687055201,0.000716566226320658,0.00212871338028942,-0.00331233255330321,0.00424613726313017,-0.00271550004147103,0.0277457514650501,0.0298003766841444
"314",0.00248689528249146,0.00166092264704254,0.0047204657733797,0.0121743617413554,0.00223173681431721,0,0.0204112087467176,-0.0018151560355405,0.00168030699048871,0.0054601548488511
"315",-0.00109455458455243,0.0054337663716264,0.000783167501147819,-0.00403308697621674,0.00911522465706316,0.00764260648105419,-0.0162881761636664,0.000909709303385853,0.00928206238608942,0.00705930535222699
"316",0.000511805440813529,0.00494716265012696,0.00704205985638584,0.0132842211406508,-0.00525178171469987,-0.00659559040390723,-0.00232379840881958,0.00999076739391747,0.0101938836565099,0.0107847322711923
"317",-0.00102235795822669,-0.00911571067161066,-0.0147628330516124,-0.0054682841278012,-0.00348400400635041,0.000110823523235659,-0.0125199576544104,-0.0151081267410563,-0.0089941868815222,0.00400083423797892
"318",-0.00723600017961079,-0.00386363835937331,-0.0149843289040039,-0.015578678643108,0.0103839716639456,0.0059753504997142,-0.0203453434473719,-0.0189917700803127,0.0214720868062444,0.0167376768781422
"319",0.00139896842206855,-0.00295549317369148,-0.00320260471997924,0.0143211846115163,-0.00335628960517309,-0.00396053934373386,-0.00210664964236462,-0.0087490282423518,-0.00563445654313077,-0.0044422060963667
"320",-0.0194091728770857,-0.0163024010083599,0.00642581322709379,-0.0163072287121062,0.00673495554712034,0.00430717230645206,-0.0036194179445278,-0.0101412848178378,-0.00512143418725408,-0.00393697157603001
"321",-0.00337392447884333,0.00197748943755438,-0.00638478578613699,-0.00236872522604659,-0.00585414888320956,-0.00252858660413913,-0.00544882337860597,-0.00986516432957951,-0.00208107331606555,0.00685105097014449
"322",0.00233236409936133,0.00488683154631242,0.00722901228883033,0.0117260727858999,-0.0124058492212594,-0.00452014205523077,0.00517433299360381,0.0136043205818777,0.00603669184461975,0.0120387266780331
"323",0.027093851038793,0.030113239939092,0.031897741195051,0.0295787065574531,-0.0097948202882443,-0.00675480880409762,0.0431490918003798,0.0302455697037949,0.0175648366762018,0.00956836643833903
"324",0.00146157757217513,-0.0128008440125161,-0.0146829021615732,-0.00725136207673771,-0.001719538474383,-0.00234050764126326,0.00580573972504594,-0.00422007683435854,-0.00761229787538231,-0.00461070342382686
"325",0.0104339821297132,0.0121388796352511,0.0274509354998465,0.0150957918756727,-0.000862663598960256,-0.00100576611871173,0.00101008999302432,0.0068176983117505,-0.0209593241348168,0.000514571753596815
"326",0.000505573021976957,0.0025442965942466,-0.00305340561352807,0.00507106371627186,0.00398925456977617,0.000111920962382328,-0.00994656473032196,0.00311169702192582,-0.00408301685887158,0.00128607698844219
"327",-0.00440280067505883,-0.00879119206717882,-0.0191424620481175,-0.00927305075392382,0.00343497561746009,0.000782849160623655,-0.00465946332358902,-0.00437875754081818,0.000221573407202191,0.00616493979980648
"328",-0.00159473952065881,0.00128032219587793,0.0109289158988919,0.0143840767823611,-0.00331690229951975,-0.00100541403763177,0.0115562224323733,0.00293175893868014,-0.0116317274276636,-0.00944611904816373
"329",0.00435674101918027,-0.00392668847173838,-0.00772199251858363,-0.0128229065981333,-0.00848104548790229,-0.00783189055651845,0.0229934864645012,-0.00877042570112285,-0.0224164982916779,-0.0167525302708712
"330",0.00925368940116389,0.00980939840410811,0.0194552974844517,0.00735355024165951,-0.00584565054609698,-0.00135301792074449,0.00339311024907674,0.00460817793402879,0.000573217145457328,0.0183485356086419
"331",0.000215099062094382,0.00072593506665708,0.01832057353501,-0.00191030237261347,0.00304908570622597,0.00180694244443069,0.00225378287585687,0.00642221553818123,0.00481270785422394,0.00231666710798772
"332",-0.00393906725723492,-0.00816452013877123,-0.00899548433525788,-0.0177044384594192,0.00379977917689267,0.001803683292533,-0.0144782894228451,0.00182300046724282,-0.0214392058059254,-0.0241397522296555
"333",-0.00589603938952987,0.0030184036529004,0.00453843020773381,0.0205983335319022,0.0071391455380132,0.00314997082969248,-0.0175439617172742,0.00873542055371668,0.00978911571586338,-0.00184207728080377
"334",0.0206857798531395,0.00729536185333846,0.00903638067253598,0.0106371423642824,0.0000651156293007826,-0.000113126897521965,0.0235192641296538,0.00739702265578979,-0.0306982566486265,-0.0232005671045774
"335",0.00276331006881914,0.00153903623180129,-0.00223867594746952,0.00958042860961039,-0.0126107259591339,-0.00810097071994875,0.00170196420285484,0.0109232603845866,0.00702469358315727,0.0253710588069842
"336",-0.00480467595039735,0.000632750113715774,0.00149567743739421,-0.000735419219841993,0,0.00147511094831176,-0.00240700554129925,0.00212603418876212,0.0199810234102384,0.0207949517827233
"337",0.00866281665284152,0.00505856043704833,0.00448099250224643,0.0111684147648503,-0.00720496041347285,-0.00317169967484998,0.00794874248949862,0.00212124669140712,0.00417294554907666,0.013151143431118
"338",-0.0178106355230063,-0.0171668331886301,-0.0126395949089187,-0.0297618312097178,0.00428870923528724,0.00397761889780179,-0.0294324498435681,-0.0225787478252779,-0.00935007535553778,0.00178157001672608
"339",-0.00258063180864476,0.00759003779083001,0.00451820183278917,0.0102929361412951,0.00897651501974073,0.00645087555149804,-0.000434840888841825,0.00721911871529235,0.0165462363085529,0.016260283314486
"340",-0.00186823120181667,-0.00599002229807466,-0.015742131921135,-0.00816391381168813,0.00369007103316576,0.00112381574766673,-0.00711326465879214,-0.00663002781526667,0.00206327377494908,0.015499896788278
"341",0.0112308444326232,0.0114132629006602,0.00380812368246186,0.0128571122150267,-0.00151392001972406,-0.00168497235660736,0.0213453219191746,0.00270573603671109,-0.00491878299974347,-0.0169866569386756
"342",0.000142539874938841,-0.004965283943831,0.00075855003838976,0.00476860642924648,-0.0109349295458859,-0.00832529502082013,0.00529622815955588,-0.00845447301910596,-0.0183929076535903,0.00550965867879594
"343",0.00206400347158953,-0.00217730475923861,0.009097853860081,0.00240625189821175,0.000437132951938146,-0.000340388063624242,0.00669195942907597,0.00598660622727598,-0.00222510835256018,-0.0161893475568939
"344",0.0125033006219664,0.0136388463196175,0.0195342162275702,0.0212723043856742,0.0090823436448757,0.00556084166451742,0.0124473518752692,0.0126241604200521,0.0211267965185493,0.0113924318653231
"345",0.000912270146785632,0.0123788380407366,0.00368455745460095,0.0127328346654247,-0.00412067716204412,-0.00169269740726319,-0.00656656267194056,0.001958744077178,0.0241379080459769,0.0145181541236565
"346",0.00273348854084676,-0.00301259078604921,-0.00146840356387712,0.00019334297118756,0.00130651082114119,0.00226144678068851,0.00759427724590478,-0.0120864702212312,0.00325478121784029,0.00148039177348736
"347",-0.00810883863983047,-0.0068432626114856,-0.00882369199086319,-0.017340213962229,0.00521977423280351,0.00304515919610937,-0.0206561727908825,-0.00791642072413823,0.0168923035786139,0.0137964968803499
"348",-0.0169147633072093,-0.00912712211369215,-0.0178040322378239,-0.010168038874469,0.000216075329261711,-0.00236166591331777,-0.0216618470915042,-0.0126952375511012,0.0116611328567406,0.0291615105691487
"349",0.000143326449162817,0.0105660104072542,0.0143505528774861,0.00291593254160594,-0.0117880790189799,-0.00653821185027503,-0.00670047066822532,0.0121234918106492,-0.0106567639262372,-0.0144037392189068
"350",-0.0134041701424611,-0.0119750577047141,-0.00819034025813714,-0.0174452711421226,0.00437720375712547,0.00442545765907854,-0.00645276198765699,-0.0098002567438279,0.00274785658118737,0.00191664407877123
"351",0.00741083861300607,-0.0038889972370898,0.00300260648001904,-0.00161416146134985,-0.00675569410493693,-0.00485756485097322,0.0143176456488736,-0.00751483052741819,-0.0204976645676532,-0.0160210091301101
"352",0.00461571500253322,0.00381346904984503,-0.0112274895851556,0.0134727678433615,-0.00888667550470401,-0.00749254601880156,0.00407460658784986,0.00757173080118823,-0.00246197401004944,0.00631828367677323
"353",0.00502484101655365,-0.00597029291994466,0.0113549774765129,0.00219331250953014,-0.00719520469175805,-0.00468997362213774,0.0104347929314863,-0.00494894936044732,-0.0295041174501247,-0.0272880294777116
"354",0.00250016951762344,0.00200231855878097,0.0134733257615052,0.00344911448205698,0.00657829895303386,0.00333353332874342,-0.00401642637843902,0.00202668219493995,0.0108657378137615,0.00670297976193712
"355",-0.0103313769349438,-0.0148943239366293,0.0022154608769771,-0.0118971089062323,0.00385732062049127,0.00594176119627465,-0.0139687329473582,-0.00845606107566987,0.00583192701538926,0.0133169815653049
"356",-0.00583156324970169,-0.00295023483134849,-0.000736726977276336,-0.0180601908724703,0.00719878650143557,0.00525609147535033,0.000729797852511371,-0.0142753371488895,-0.0122783311991624,-0.023606741866913
"357",-0.000506784779923164,-0.00989353350327737,0.0117994298243056,-0.00871917956155954,-0.00890585388742349,-0.0036370446977827,0.00554624812219684,0.00921574779590206,-0.00264727219085892,-0.0149551263085738
"358",0.0199970766244697,0.0193311696853109,0.00801739750844876,0.0318166900430308,-0.00599091196732371,-0.00524769552911875,0.0251089441553751,0.00913152031209297,-0.0023081938301629,0.0379554310072467
"359",-0.0318936547009288,-0.0281265297071146,-0.0354302945210627,-0.036230412070832,0.0129464578658638,0.00871584707174522,-0.0396430669136157,-0.023268833203281,0.0301908743848771,0.0255972879346751
"360",0.0024210402872149,-0.0010367562313407,0.00149913294109671,-0.00255696292092511,0,-0.0071628805557129,-0.0231462825262843,-0.0138019950188428,-0.0120143726030624,0.0102211742407385
"361",-0.00497722660539557,-0.0136831995423764,-0.0217065804282153,-0.0230703028485716,-0.0065005618358932,-0.00595397181973356,0.00392404104995236,-0.0279905751162335,-0.0277303677174762,-0.00400007566573857
"362",-0.0147122407599711,-0.0154995568800953,-0.0145370454972829,-0.0149637939618114,-0.00232967969235254,0.00103683087993978,-0.0205953438446403,-0.00394509718179681,0.017182863219771,0.0368531702795376
"363",0.00380751654039968,-0.000874282014111993,-0.00232915245800769,0.00583166993565376,-0.0100041789099649,-0.0087458114831872,0.00613981210664694,-0.0128711167336001,-0.0163180768668609,-0.000227787839221172
"364",0.0126440056810198,0.00787874748349116,0.0101166045131891,0.0108082238012779,-0.00213352364802877,-0.00232182835021788,0.020899626313446,0.00902712645860992,0.00268696267960178,-0.00638108513231939
"365",0.000587998942909174,0.00550080302791089,0.0092451633103916,0.00339914365454952,0.000224816061243027,0.000116226748140713,0.0143456564055198,0.0069582287762513,0.0137481064022347,-0.000917259715971785
"366",-0.0048450887105348,0.00124744182106307,0.00687006356730047,0.0042338585455941,0.00202465511698779,0.00337393430451072,-0.0294636485484476,0.00592292736706757,0.0027582805939943,0.0101008964033154
"367",-0.00973624581991195,-0.0107360626962452,-0.010614081811999,-0.004848954848648,0.00842109972572214,0.00544957124837619,-0.0148754972672005,-0.0107951224702459,0.0118051461318052,0.0136363564003168
"368",0.00126584503335403,-0.00164741979216065,-0.00306482414856324,0.00155391111794345,-0.00590043058253131,-0.00576589499478319,0.0206465816925456,-0.00297607663388588,0.00158585185303406,-0.0233182687419895
"369",-0.0162314219003633,-0.0197998005331145,-0.0330517196943719,-0.0326449124131449,0.00582400839750497,0.00464048949178597,-0.0247578159403912,-0.0107121542683088,0.00599410780353082,0.00688701191158803
"370",-0.000988136137223705,-0.00372102759825332,0.00715394411003478,0.00291535026883305,0.00211527256027044,-0.000462186918460006,-0.0207429255105516,-0.0207612264464411,-0.0209106358935571,0.00706784901461277
"371",-0.00197807974173059,-0.00377547908888631,-0.00789257411615407,-0.00443308579577373,0.00666546077728558,0.00531376844084663,0.000473852126449792,-0.0022866603377284,0.00436335994320181,0.000226438523680317
"372",0.00472589895284381,0.013418223833263,0.0151879230033283,0.0200241479330237,0.000442492767840585,-0.000116301523400142,0.0176522265854895,0.0177083408968977,-0.000571658847928758,-0.00384796818793998
"373",-0.0271600478193186,-0.0245604580280061,-0.0251966049302363,-0.0343104808988878,0.006729722732145,0.00563231794482721,-0.0357588771710552,-0.0227228009415239,0.0364905407570473,0.0331744203459301
"374",-0.00545895528367524,0.00466262676213614,0.00565392542695919,0.00966896586276222,0.0117260520110138,0.00491330557549063,-0.00780687353263243,-0.00691238024990404,0.00949122602923258,0.00263902291314744
"375",0.00352849683373013,0.00268149039453958,0.00160673668523104,0.00757294191785607,0.000217131995107422,0.000681682379875204,-0.00327911143199588,-0.0101242841182188,-0.000765267292388017,-0.0177670229074153
"376",0.00312566687840699,-0.00874319717259509,0.00400969133837847,-0.0178312105233003,-0.00236997296697938,-0.00271332313236905,0.00575668010998909,-0.0100149385494493,0.0137855795670552,0.0176417854465454
"377",-0.0171367769563691,-0.0153574116380706,-0.0215656326218261,-0.0285067936005825,0.00522985239730356,0.00240110084288125,-0.0207684371891301,-0.0079636807646134,0.00550392810257172,0.0190915051542797
"378",0.00103042458738689,0.00779865157709891,0.00326519324393604,-0.0028573862705451,-0.00216771623713741,0.000342398251591769,-0.00801629660297443,-0.00282072284157864,-0.0119137063843235,-0.000430672741844051
"379",-0.0102128583453489,-0.0119209760412033,0,-0.00356240004459984,0.00456166496642507,0.00467461716104656,-0.0205383957005767,-0.000217683188597384,-0.00901580510570943,-0.013571687391414
"380",0.0177570767533823,0.00910145629617376,-0.00406812152626612,0.0122795497007875,0.00648720089380372,0.00249627293837551,0.072361252901586,-0.00217604168830665,-0.00405570522671139,-0.0362524577358925
"381",-0.0192552026271411,-0.0098585506669262,-0.0163398239260212,-0.0201919350233253,0.00440444785021521,0.00475468115356836,-0.0735694749468707,-0.00719723112665738,0.00704379257050647,-0.000679765429519197
"382",0.00408711664585715,0.00646132803154997,0.0091359331813512,0.0181009787542414,-0.000107101913953023,0.000337304629694613,0.0181661243504623,0.00395391639049003,0.0221857814207651,0.0272107961405996
"383",-0.0116520792395284,-0.0181014719097066,-0.0131687958148707,-0.00669606493114849,-0.0142261950856514,-0.00934755296477707,0.000340045074035844,-0.0205687226562405,0.0174276169937733,0.0139072576091852
"384",-0.00904405510515527,-0.00321538434047608,0.00667240298333427,-0.00123972966769981,0.00878973644581249,0.00534348067722501,-0.0348223067762514,-0.00379792257377121,0.00788146246820243,0.000435523166912199
"385",-0.0140971261289644,-0.0148385225772862,-0.0165700399495838,-0.0166799304574792,-0.000323368727587203,0.00361810398620466,-0.00950395019931494,-0.0222026428657347,0.00271081210673296,-0.0317736170793276
"386",0.0245475569516675,0.0128791046342103,0.0252736693947904,0.0288759856893639,-0.0180758896396299,-0.00912637284886331,0.0701849088095166,0.0155964541340976,-0.0179889366328155,-0.015284340931413
"387",0.0100032203255931,0.0223062631444926,-0.00493018630361519,0.00467739122628941,-0.00514995765911364,-0.00477608191028167,0.0161046782881622,0.0219058089178112,-0.00232953192864194,-0.0235107378302527
"388",0.00623006450956676,0.00980250382840131,-0.00412858943541428,-0.00862460410232413,-0.00374557677140752,-0.00342751210084236,0.000326799277783119,0.00773499292244129,-0.000530704727969455,-0.0170640232062798
"389",0.000555471017086751,0.00584576506424805,0,0.0123954169120324,0.00387073709718222,0.00229303432546857,0.00294020571263642,0.0164471913093296,0.0100881917826949,0.0121285500252375
"390",0.011344784139218,-0.000104047860824963,0.0132673456837005,0.000608171693123882,-0.00495690868970888,-0.00343178123148258,0.0317590478440652,0.00539390891588676,-0.0216569063817208,-0.0218516034181685
"391",0.00541274400577363,0.00352906075627613,0.00654631663253347,0.00144378001780443,-0.00199133256560513,-0.00160588925311667,0.0213102642002803,0.0313304269854897,-0.0267569100957857,-0.0225799169704837
"392",-0.0207537194555674,-0.0212017841325874,-0.000813165287574136,-0.0369581416057291,0.00975813772723577,0.00862166173891254,-0.0615148001971851,-0.00728249617207444,0.00839132162967871,0.000737439518115224
"393",-0.000239228141538983,0.00612835282109758,-0.0113913782201995,0.00685533885295442,-0.00999389865855715,-0.00581329048012114,0.0151515751955504,-0.0253613140873827,0.00394174961257554,-0.0125246920014604
"394",-0.0146636824467536,-0.0149127814274925,-0.0115224618549152,-0.0169049255766658,0.0100947849159874,0.00573266952827534,-0.0212527550573254,-0.01096762757253,0.000436263487048283,0.00497402307860817
"395",0.0213525068760547,0.0110872437715743,0.00582828709709204,0.0554092681265497,-0.00406387435071331,-0.00285045826443431,0.0500583431113673,0.00217423237812708,-0.0124278530765991,-0.0113834159100783
"396",0.0178174470840353,0.00991147525022162,0.00910616237044137,-0.0104094178015316,0.000993103201280654,0.00194441465891337,-0.00489322988164154,0.0197439256027891,-0.0118114477011346,0.0197747231077408
"397",-0.0132263604992983,-0.0110668621573836,-0.0155866172112846,-0.0224103329137525,0.00991549005527381,0.00798664768293067,-0.011739009148139,-0.00531931043827449,0.00625564140713708,-0.00834558517007378
"398",-0.00528287168102259,-0.0130911800238789,-0.0141665948093299,-0.00678378276532032,0.00221102542688634,0.000499766669858071,0.00240786442414853,-0.00342241857290793,-0.00566165617980341,-0.0111386394825681
"399",-0.00927379849213561,-0.00363731611973861,-0.0253594308856314,-0.0306164293878493,-0.00229436475250178,-0.000680932912637044,-0.0140911167542096,-0.0223224072682821,-0.0159651780730155,-0.0330412197272842
"400",0.026961934594335,0.0300622495478773,0.0225500416445392,0.012876296822445,-0.00744498317202291,-0.00511274635611447,0.0427154328884021,0.0208564385968686,-0.0233718745560686,-0.00698947251736459
"401",0.00444104632005815,0.00145939834408515,-0.00593722265845387,0.0199089843331641,-0.00408187404827731,0.000342101825330232,-0.00467284717208194,0.00559157877414496,0.00650554120572644,-0.0106882484373897
"402",-0.0148920355802404,-0.0185264395910536,-0.0221841800759009,-0.0343370761193377,0.0162834843092736,0.00936116269889098,-0.0242568285973189,-0.0248079629295906,-0.00634814180918908,0.00553359520466379
"403",0.0185814861095384,0.000424370451486356,0.0148340216998675,0.00243591336832738,0.00272381304352698,-0.000452065076902319,0.0323980517484783,0.00197372410256746,-0.0192821010236776,-0.0280398631922217
"404",0.010357599710844,-0.00190788363677019,0.00601861698930906,-0.0104475257975186,-0.00956503181526414,-0.00486601778944784,0.0245451192251345,0.00656633252370664,-0.0390856686012081,-0.00107836893611957
"405",-0.0104046590395537,-0.00488547303167808,-0.00683758019810266,-0.00834757323165758,0.00932913640334099,0.00693654835086854,-0.0221377681659183,-0.00478405222738409,-0.00751879727050897,-0.00863694178083629
"406",-0.00603011256365116,-0.0175027606361129,-0.0172115579827478,-0.000247587341732025,-0.00347978377180158,-0.00214490330830031,-0.0161266258305396,-0.0190080454938174,0.0129160586034298,0.0334875668411299
"407",0.00754457235742567,-0.00695183518723907,-0.00612929283338826,0.0131250271520043,0.00643728379407515,0.00305436423403527,0.0165488087736789,-0.0144764183357673,-0.0270966166526879,-0.00869334665424149
"408",0.00486324562276508,-0.0070006270726779,-0.0070486414898846,-0.0156437103807896,0.00867335732449925,0.00372351543415439,-0.00155044741741783,-0.00338998581073546,-0.0216761316112446,-0.0135530788405448
"409",-0.0136742414750942,-0.00638937553388363,0.00887305029385788,-0.0168859782963803,0.00397678806721169,0.00247228727145687,-0.0209625065240795,-0.00680294599674813,0.0150715708516644,0.00565732592459312
"410",-0.0109042328942185,-0.0121949888809805,-0.0158311493739985,-0.00833574175023744,-0.00385363760321833,-0.00145717618106422,-0.0206186167963465,-0.022830911349251,0.0206852403292421,0.0155371930081818
"411",0.00464583016929709,0.00224484905947175,0.0107238164683165,0.0254712899484284,0.00279378744641945,0.00291951144349145,0.00242850927036198,0.0163553052918237,-0.00460029839612097,0.00791332262534139
"412",0.0017243072897235,0.00515100347219821,0.00618933567180946,-0.00148996825990233,-0.00182153901918869,-0.00212810399229379,-0.0137314440323307,-0.0114945132943785,0.0279790788903094,0.0429208050077479
"413",0.0144756188005914,0.00713009594271474,-0.0070300611353088,-0.000746754047422304,-0.00064496838342909,-0.00291643415694187,0.0229320201240359,0.0090700419653349,-0.0148238269201523,-0.0338770128588113
"414",-0.0202849970155842,-0.0163716751938718,-0.00884957584739499,-0.0206620743090962,0.00999188393886707,0.00663781479656356,-0.022097884742413,0.00230473961868682,-0.00185004928835575,-0.00571443886543999
"415",0.00291282401348836,0.00382387828595476,0.00535728428814575,0.00177969712697634,0.000850920322423399,0.000336678791056588,0.00769609198207766,-0.00436896718114477,0.00370694427282814,0.000522586882356402
"416",0.00973341533609506,0.0109790572070287,0.00444043851715459,0.0213141671846959,0.00170051526922088,0.00145183223356748,0.00893777183918276,0.00808342302194798,0.00160036926257412,0.00939941240979691
"417",0.012128348691121,0.0141843703260029,0.00795740637787112,0.00695652625685783,0.000105637357445731,-0.00144972747249295,0.0331770043406001,0.0119127074527881,0.0100786503186008,-0.0196584834087645
"418",-0.0107536205508914,-0.00611883247105494,0.000877282844706118,-0.0118433962262949,-0.00445539072467016,-0.00122930813825994,-0.01122342895644,0.00271665536991827,-0.00571916524701888,-0.00369406808285622
"419",-0.00621178612265305,-0.0127530538263563,-0.0131462435600133,-0.0302118874788641,0.00930461256412163,0.00544398552020331,0.0122971180531231,-0.00541898375988015,-0.0307184191741331,-0.0259532462648115
"420",-0.000859507902782219,-0.00467672007889408,0.00444043851715459,-0.0164777776843518,0.00423902732200743,0.00245627827034278,0.0137048009771457,-0.00726420998991073,-0.00391411630987804,-0.00570970809837212
"421",-0.0301061015735163,-0.0449767508428891,-0.0318302435019444,-0.0460732985354702,0.00801959225439552,0.00501123475677168,-0.0311875318441525,-0.0420764419771621,-0.00633793898260793,-0.0142191914588167
"422",0.00314438036983855,-0.00562310234750873,0,0.0142698228401119,-0.000524081208020055,-0.00221631295058378,0.0063432549787934,0.00501309214160872,0.00752652133596787,-0.00998620532375682
"423",0.0206559780421156,0.0172008743202503,0.0246576976442885,0.0124460587259509,0.00418964272780209,0.000110510414742304,0.0431770554697104,0.0261284571030778,-0.00151939725806294,-0.00224151519185878
"424",-0.0296875659721261,-0.0277972442246801,-0.0276293740767004,-0.0561199089699985,0.00990800860576657,0.00455389952567931,-0.0438067912400708,-0.0199073431015574,-0.0300532966008965,-0.0365066424621719
"425",0.00405791478847184,0.00428887534243327,0.012832183759746,0.0161382885922021,-0.00619617670528894,-0.00254266323343744,0.00537138293993134,0.0243269671110884,-0.0296770435266582,0.00145725716199618
"426",0.0144680785358977,0.00142328154063098,-0.00542959501376017,-0.014767278343633,-0.000519588355200717,-0.00177324063869799,0.0114707466230464,-0.00807024010396307,-0.0153597276292141,-0.00844003600158705
"427",0.0046209740573524,0.0234543883983578,0.00636955162367148,0.0333708486579725,-0.0128931562920354,-0.0049963163516582,0.0105638074370527,0.0167364218239567,0.0337985896606847,0.00675078805886775
"428",-0.0475848299944177,-0.046759288811672,-0.0280292907089424,-0.0785441297900131,0.0324423056500054,0.0191924198235716,-0.0614911841514757,-0.0477824947542697,0.026604830181145,-0.0393584528508193
"429",0.0167372726394794,-0.0118991106100664,-0.00930234464643165,0.00861305550178693,-0.000204388613479711,-0.00284649489423505,0.0307943923139524,-0.0177671241212914,-0.00992775941020507,-0.020333922337049
"430",-0.044963062226579,-0.0459569109377364,-0.0356806937300451,-0.07096580708945,0.00500043609299161,0.00900336036908334,-0.046559769335505,-0.0381325454457248,0.11290529869898,0.0300495994542949
"431",0.0296714739964827,0.0569292556894478,0.0447905589189774,0.084310660808798,-0.0146211147861154,-0.0117519566602207,0.0845001556800844,0.0200763663933543,-0.0311256263880836,0.0018046140202741
"432",0.0397139958478068,0.071410785011139,0.0540541505003778,0.124525164677874,-0.0317357323448022,-0.0178378516192256,0.0327337748200114,0.0652989271150723,0.0384057957099349,0.0330228692629901
"433",-0.0226395868914858,-0.0204729750723708,-0.0344826585562673,-0.0652458824419585,-0.000106371417559092,-0.00212980367941473,-0.0880947575643575,-0.0179792483670932,0.0372179214741364,0.0345829335306627
"434",-0.0227515181195052,-0.0234552782247822,-0.00915763790375079,-0.0311454914252647,-0.00383211249585313,0,0.00636368609519633,-0.0158998080893874,-0.00964341780668332,-0.00983125370641769
"435",0.00320522983004756,-0.0019028467568778,0.0138633989287509,0.0114810787595356,0.00438070743299201,0.00258406897993102,-0.00739023031371855,-0.00612064515083111,-0.0182291779891304,-0.00822696864585204
"436",0.0156396710027655,0.0243032167180401,0.0173198211132,0.0513618409945653,-0.00202148519159018,-0.0030257623554929,0.0185308243030757,0.0187197375565189,-0.00299852384959665,0.0174484640515546
"437",0.000496480017237122,-0.00930453308428236,-0.00537637658669554,-0.0340079324155962,0.00724799854718539,-0.000674149060217566,0.0207926907539309,0.00580240269627108,0.00219782540883151,-0.0118076703580804
"438",-0.0783614838586015,-0.10354549000007,-0.0774776015887485,-0.116792505963998,0.0291006970609902,0.0139463955567802,-0.0598344220211082,-0.0973555490220709,0.0338181098086114,-0.0620198269049511
"439",0.041389882025715,0.0440024193134718,0.0410161468938453,0.0809869317942369,-0.0243695334864982,-0.0132004971082953,0.0485781616199448,0.0162449283182604,-0.0502400357262476,0.0279040396033075
"440",0.000603292687778811,-0.00125492242276493,-0.0121955099313872,0.0119990457609744,0.0125803931287674,0.00704968814607954,-0.0153347643846783,0.00943414444230495,0.0105795345009991,-0.0233106248146986
"441",-0.0362741147389916,-0.0419491768693858,-0.0427350871342106,-0.0876230253731889,0.00803922721911121,0.00560078846365575,-0.0662297511573826,-0.0501041215787444,-0.0423403391608662,-0.0552870733393158
"442",-0.0135002109198202,0.00209792193288227,-0.0198412210304988,-0.0263073030982273,0.00880341653361083,0.00378754546456794,-0.0533708044125939,-0.0213173477157439,0.00315794963784888,-0.023345023034933
"443",-0.0509336894390425,-0.0580848772094748,-0.0323885642216831,-0.0751953681425761,0.0181721378530495,0.00809931588097479,-0.018360242206568,-0.0823790818693318,0.0204625630445605,-0.0425672076916122
"444",-0.0447859913123761,-0.0500000139489841,-0.03661090220258,-0.0777895118071785,-0.00302430920411334,-0.000769616361279812,-0.0844511580144839,-0.001826138199711,0.0354769581807897,0.0123118879564208
"445",-0.0251924245090427,-0.0102343173457277,-0.0369162435714957,0,-0.0143629730819668,-0.0127787953076347,-0.0167152385192101,-0.0423780788829878,0.0246361988530834,0.014527083835969
"446",-0.0698393279924893,-0.0747412347278782,-0.0462232156224829,-0.0736640177901864,-0.00841455237018185,-0.010041369993925,-0.0715631405424936,-0.0799106929849241,0.00536797149111989,-0.0466200320130208
"447",-0.024255353293509,-0.0249042307067888,-0.0437351992803768,0.0115367235773118,-0.00703734403011147,-0.0117235095115643,0.0795659331764678,-0.0311418098450797,-0.074304792562741,-0.0443590389076348
"448",0.145197548316608,0.137524678312813,0.158219794975282,0.227698626789179,-0.0128189868635205,-0.0068423294449701,0.0747486168894751,0.107143081748968,-0.0147801368086982,0.0555555194676047
"449",-0.0148001004476587,-0.0184227780909215,-0.00533607632239941,-0.0497676272150791,-0.00644040502185528,-0.00470873095967927,-0.0648743130662957,0.0438709627228235,0.00256127582781485,-0.0183518618979334
"450",-0.0984476651138143,-0.105571734978651,-0.104077255632865,-0.161662120671408,0.00956399633042104,0.00819233546591347,-0.14166664519549,-0.0908531636396415,0.0135036622933209,-0.0455026021484503
"451",0.0416572179015977,0.0498360218641278,0.0610778969192574,0.0491461254510577,-0.00515778507976605,0.00022854723903154,0.062864155322381,0.047246928907658,-0.0482534761314001,-0.0188469788539656
"452",-0.00597190844268047,-0.0162399509047457,-0.0135439261556817,-0.031361511123806,-0.00687711729781848,0.00629288237796133,-0.0102767075145079,-0.0327815538009583,-0.0262328411371821,0.0112994087772322
"453",0.0600795161035814,0.0520634527044823,0.0789470079108063,0.0700818544260251,0.00799026558399141,0.00102344856220316,0.00946035784903687,0.0620804900339498,0.0167076935203692,0.0201117479402557
"454",-0.0298554662731325,-0.0585395711525618,-0.0360549018248038,-0.0796630891601503,0.00528389799494566,0.0105638921884157,-0.0345141911152462,-0.0423380226274573,-0.0314649808917197,-0.0357795082209367
"455",-0.05445385017813,-0.0762819163022954,-0.0605060768645876,-0.105285148104259,0.0202911506763244,0.00764270821701807,-0.0733899671541098,-0.0514680790064955,-0.0568196771908416,-0.0473305935845669
"456",0.0115837112529051,0.0183901275456537,0.0339577905984108,0.0279073110054675,0.00741839690985735,0.00133965450478435,-0.0155854266936972,-0.0285219746789565,-0.0147817182370898,0.00397460927152582
"457",-0.0507142685087612,-0.0494037930072643,-0.0600224506953867,-0.103167723481773,-0.0106374547129399,-0.0042341459307268,-0.0641056970246578,-0.0748298527207426,0.022080636317604,-0.0399841171555951
"458",-0.0355005969073288,-0.0580646017264962,-0.0602412483800925,-0.0262358795996136,0.000723947099786404,-0.000559336374910901,-0.0521354332250806,-0.0170280197192976,-0.000415441080396484,-0.00742275787031688
"459",0.116854954256817,0.129756536397139,0.1217948995166,0.209326393889737,-0.0145665002292269,-0.00805937508365773,0.163253477616466,0.0362206249324153,0.0223053615960098,0.0274200670797233
"460",-0.00725272179126701,0.0148198036877256,-0.0228570487876592,-0.0317051188840335,-0.00503186496559438,0.00146722520852638,-0.0397387169751087,0.0136780030800543,0.00284590048995925,0.059037684233568
"461",0.0345940790819856,0.0288749613573858,0.0538009074476733,0.134956110958515,-0.00906064084125613,-0.0076616557525101,0.048454867735205,0.0468512987598091,-0.017432445945946,-0.0412371829495353
"462",0.00550338954643159,0.0125805602107882,-0.00110968801041145,-0.00857764381566317,-0.012972442978332,-0.00204421119054232,0.0629527587735403,0.0204081478810851,-0.0188420164879936,0.0111509323669647
"463",0.00289159933787109,-0.00382300625111642,0.00666650391665335,-0.00904407966655896,0.00270391998197894,0.00159826251617723,-0.036427682825375,0.0245614996523509,-0.00336414372661309,-0.0110279603272104
"464",0.0339824719104687,0.0697156018408336,0.0551877866495505,0.0912698524495452,0.0187682879744713,0.0119721627310221,0.0556096309482776,0.0352737580864686,0.0616034475837819,0.0454003257497158
"465",-0.0420276768956299,-0.059491884768034,-0.0209206063662299,-0.127272774211961,0.0118579745755618,0.00529425033014386,-0.0965801130199091,-0.0370491467601426,-0.0355060929184117,-0.0259048539988933
"466",-0.0554115140067435,-0.0632549555071528,-0.0865382917116441,-0.0504166607727773,-0.00721967192031214,-0.00302545261943032,-0.045268844972437,-0.0398483500573027,-0.00796706011124759,-0.0438013163797875
"467",0.0330181679096802,0.0563286847239119,0.0584796768287499,0.0811758676038798,-0.00653456466748847,-0.00359733560851394,0.0592020772111093,0.0296949160249347,0.00387702847027116,0.00122699958366002
"468",-0.0131046637754417,-0.0215226731254043,0.00883974056591086,0.00933425542395749,0.00488073522768984,0.00101562495499397,-0.0857363485943994,-0.0535088668463697,0.0148965793103448,0.00653592119552315
"469",-0.0308757315117446,-0.0252791562033579,-0.0416212163029904,-0.0623239577708339,0.00295536217742542,0.00371877801840292,-0.0127245935208671,-0.0326726541377507,-0.0207936797827213,-0.0190745666179768
"470",-0.0440011645288737,-0.0565846918101029,-0.0274285974663695,-0.0741852001017608,0.00642058227819087,0.00617620053780077,-0.0736901666865765,-0.0288422886190112,-0.0284525040200208,-0.0293754072624588
"471",0.0623394234944186,0.0828274988595226,0.0681552971898631,0.138489993085485,-0.0239502431446501,-0.00725393668817942,0.110708046084282,0.044157722414307,0.0307143142857143,0.0187553871036426
"472",-0.0499059858149423,-0.0524234505141269,-0.0539053780712953,-0.0960130028187652,0.0198237566380608,0.00989218722658869,-0.0985837533987162,-0.0550149569772006,0.0159390293571995,-0.00627609242624128
"473",-0.013276965786133,-0.0327068294697089,-0.0023256421240484,-0.0166513465432824,0.00441304981347446,0.00422978812584218,-0.00785528162370197,-0.0213863993173454,-0.0088676804010499,-0.0227369028419511
"474",0.0188370569461687,0.0143884546783264,0,-0.0146454997548017,0.0128677642624617,0.00775895147531513,-0.0401947871147434,-0.0129499851238185,-0.00192704743490579,-0.0150796573222827
"475",-0.0640789430073369,-0.060638099719699,-0.0641025949801616,-0.0863912878341623,0.0256142923559337,0.0107779601782807,-0.120558474040661,-0.0873311466723421,-0.00344780020830782,-0.0113736460813515
"476",-0.0742331359346956,-0.0683278562868648,-0.0286426786527263,-0.0716826263773958,0.0516615520645234,0.0201312666740809,-0.0873018370287436,-0.0336921791110484,0.016468239234203,-0.050884855047417
"477",0.0539429473894837,0.0571314744602658,0.0615383656362649,0.144030290511459,-0.0144597022637665,-0.00917376353348687,0.0826091358229879,0.0418406441548014,0.0735194175705685,0.0172494312916369
"478",0.0692909760403564,0.0770406042128604,0.0471016829162851,0.0607947913024174,-0.0156432732990519,-0.00936613575894407,0.14457812428056,0.0441767092283893,0.0261256316074987,0.0687441540990277
"479",0.00740918051125661,0.0202850093675084,-0.0046139411713737,-0.018953171266304,0.0294151606037516,0.0171706368569753,0.0271133388046934,0.020940113368118,-0.000494388802650403,-0.0334477063449429
"480",0.0386406011202298,0.0177884811228683,0.0185402568171045,0.0763575454885246,0.0013422473352136,0.00609049628604708,0.0456521816034459,0.0397658580076123,-0.00605918117747561,0.0319432230558587
"481",0.0125888743601326,0.00342723032164849,-0.0147894546621956,-0.0192310301971163,0.0123528079173536,0.00201653616662156,-0.00861303301512029,0.0362318086785434,-0.000870850990452365,-0.0434221329352545
"482",-0.0885777988647102,-0.0877732914537159,-0.0577368614054388,-0.0962962937965063,0.0382953633350251,0.0135359902611802,-0.206111723687275,-0.0784771274728431,-0.0580251041719612,-0.0310112387636797
"483",0.0384843729359494,0.0490449064695422,0.050244985310862,0.0631626779386618,0.00383940896328938,0.00524548555604243,0.137735890998853,0.0408939316547603,0.017184335302463,0.000463807880641598
"484",0.0240415165019103,0.00749471658017087,0.00933499374826741,0.00816342730941799,0.00282182738135828,0.00156533342329168,0.0454398647649414,-0.0064805063469735,-0.0100064591295564,-0.0115902577741106
"485",-0.0231333036829957,-0.0262130359848585,-0.0393060921108763,-0.042734980697662,0.0197050029337185,0.00625164312063076,-0.0164974172465174,-0.0342438197670699,-0.00892622735626158,-0.052532722436711
"486",0.0308318851783982,0.0152783167306845,0.015643423445556,0.0592108387907966,-0.0162066015593975,-0.0105620014026525,0.0964515178905463,0.00253284399542508,-0.0129801721854305,-0.0247524516760373
"487",0.0349144672227175,0.0458616070701079,0.045023768779662,0.0638859979505948,-0.00217256776241925,-0.0037671050464344,0.0941450673438693,0.0484211230425975,0.0225442843214285,0.0461928228227908
"488",-0.0164833096728879,-0.00548140481132264,-0.0068025556123178,-0.0137614881376672,0.0197752503603241,0.00850999058261204,-0.0717931785458219,-0.000803433208772519,0.00170610242937408,-0.0218341123036047
"489",0.00681519197509206,0.0285912218224003,0.0216891804321455,0.0596195541470386,-0.00240154883960209,-0.000938481982047046,0.0663381887387455,0.0478292514823961,0.0448054226436416,0.0302580101527612
"490",-0.0240811355162314,-0.000669951734933893,-0.00335151773429843,-0.0255385850504168,0.00196140726805671,0.00604690033700828,-0.144254216794447,-0.00460234832389383,0.0112852915360502,0.0317765472120874
"491",0.0119394683505505,0.00502692469912014,0.0224211202734628,0.0139231389069374,0,0.0027987585489333,0.09460320156476,0.00346805281583551,0.00198383132092173,0.0219319417556862
"492",-0.0139338329937352,-0.00200085597195432,-0.00548241774049218,-0.0133282763708212,0.0113906077587818,0.00217007149027726,-0.0284225291942174,0.0145929688930451,0.0221507244685244,-0.0282931297013179
"493",0.0470654217219839,0.0648181504281897,0.0507168807941616,0.0798201124083453,0.0247249832755303,0.0158813405381428,0.121791106547144,0.0264948865507211,0.0225181724580672,0.0143198584309669
"494",-0.00968657021970754,-0.0097270570662028,-0.0020987545705875,-0.0174374451960415,0.0271341085834365,0.00680105230671679,0.0252794516649579,-0.00921813799145765,0.0114847384736532,-0.0136472101417828
"495",-0.0186830653343337,-0.0323193549030883,-0.034700348722655,-0.0219908048358277,0.0209827801878306,0.00675541307373351,-0.0788995435818746,0.00446553420223506,-0.0182605290881425,-0.015267213431192
"496",-0.00430226732573857,-0.0216110235622686,-0.00435714831921963,0.00355031447853915,0.00106493541951669,-0.00330482926586628,0.0495913779802402,-0.00156732464611442,-0.0147848569887377,-0.00678285373721177
"497",-0.0128128108188357,-0.000576061926008897,-0.00218844055465195,-0.037342810237228,-0.00768892290433909,-0.00261221125232436,-0.0209396541243355,-0.0332709756759678,0.0100448024946678,-0.0282925977976181
"498",-0.010337658314141,-0.00576470836372778,-0.0171363040836534,-0.00828138787368093,-0.00131887665253538,-0.000503926935774279,-0.00759253028166218,0.022814758170411,-0.0099449078593925,0.00401600906206068
"499",0.00580294389763125,0.0133013574094747,0.0123733022264418,0.00709809618677149,-0.00214559630131461,-0.00100816470695075,0.00765061782920395,-0.00189029629703064,0.0100448024946678,-0.0154999422095188
"500",0.00576980188017107,0.00807824443134586,0.0188893795236695,-0.00331657971100763,0.00330824281199926,0.00534788184791379,0.0132175439744084,-0.00378732075196853,0.0256410139664631,0.0157439728792961
"501",-0.0028682927014505,0.000333844973501973,0.00763294524796332,-0.00166425807876802,-0.00119888810961677,0.00220637354542585,-0.0563422334759544,0.0112015040428302,0.00876168244770281,0.0110000038080995
"502",0.0237025406689224,0.0283711830317885,0.028138703160643,0.0266665789774325,0.00952332993069827,0.00140647957575446,0.0452942138913162,0.0113036081756854,-0.00521130295799199,0.00593463684071205
"503",0.0142745985209252,0.0107107955071426,0.0084209595927629,0.0133929692271306,-0.0209185039215972,-0.011040378630323,0.0475520205210069,0.0089417976746875,0.00721763661891428,0.0417896661742048
"504",0.0301418150578165,0.010597290099952,0.00521925567742976,0.0476571326674686,-0.0251364353325576,-0.0143106843571337,-0.0273972304994362,0.0347118605047498,-0.00335175693545164,0.0349221404623925
"505",-0.00118341994409665,-0.00953282421549939,-0.0249217815219395,0.012996850865804,-0.025784205271049,-0.00175057752846797,-0.0196079823269319,-0.0071380908109151,-0.0202945603515751,0.0104879131647666
"506",0.00667739014812452,0.0121912083588338,-0.00958506528788194,0.0226417738943878,-0.0100572257573145,-0.000618598334330644,0.0495777450726944,0.0273187336443235,0.00769405749192509,0.0261732517063458
"507",-0.0299558946994034,-0.01172750316982,-0.00967714733976721,-0.0575645661476069,0.00392080891561575,0.000206192890617851,-0.033816783897236,-0.0129457741418092,-0.0279572076103797,-0.0510114152463199
"508",0.00408088963042941,0.0128288319728374,0.0141149789106514,-0.00430705432780509,-0.000798625639203521,0.00268316141635427,-0.00444412945801298,0,0.0206646404833837,0.0037070854943253
"509",-0.0214195577314993,-0.0345158598411773,-0.0171307533770876,-0.0216279759483929,0.00151055134113154,0.00463094880910098,-0.0460380779579366,-0.0212692980783469,-0.00639357099684534,-0.0115419980752803
"510",-0.0240207349311748,-0.0272215064948004,-0.0119823613369034,-0.042202787975766,0.0103788093073682,0.00624911407466011,-0.0582039624989136,-0.0315100881933605,-0.0376548626705163,-0.0453058901349086
"511",0.00184012211710183,-0.0188807348547652,-0.0187431944045092,0.00293762476358639,0.00105301596496665,0.000712121381177377,0.0301239496467065,-0.0373973281129588,0.00148582215240656,0.0166340748254159
"512",-0.0314539796735626,-0.0474230244459817,-0.0292133536251865,-0.0485353513242666,0.0164888361262077,0.0055949762491363,-0.0518538959985972,-0.0470087229818827,-0.0134767067313318,-0.0139557828393829
"513",0.000355116015327894,0.00649365817196523,0.012731360278474,0.0114333329582901,0.00163900535829287,-0.000809102170561848,0.0289348258967759,0.00163096426626863,0.00751971415566222,-0.000976072559683128
"514",0.00782024645738555,0.00143365167601539,0.00685748860302948,0.0108695297251475,-0.0154186629873238,-0.00921329999194265,0.0367735792845247,0.00488399960735375,0.0288593112185509,0.00439661793669699
"515",-0.0527863097048781,-0.0776664024327907,-0.0431330364627536,-0.0744085260438957,-0.000174945821604044,-0.001533004828566,-0.108196371187102,-0.0810042145617409,0.0218836660849193,-0.0311282811770387
"516",0.0431921163661129,0.036476355993101,0.0438908877540032,0.054368145401134,-0.0315894040093251,-0.00890394052782639,0.0995985030437088,0.0599383022351483,-0.00437760308959789,0.00401600906206068
"517",-0.0154668945057863,-0.0243352694552776,-0.0249999674634781,-0.0330543762876694,-0.0192468586109438,-0.00660868363207967,-0.0507599884485459,0.0112262019820739,0.00510992263553356,-0.0129999764309525
"518",0.00435034123728917,-0.00652334737363025,-0.00233093215858782,0.0127620949494434,-0.00783071909482458,0.000208280033457742,0.0317004293297294,-0.0143911220469064,0.0467013112626791,0.0466058108368732
"519",0.00685845876760038,0.0266513041325884,-0.00116831228097891,0.0117013610551597,-0.00872881872025766,-0.00249405662083346,-0.00838008112284905,0.00709187319457971,0.004744131986266,0.00193618162824372
"520",0.0101578482999116,0.0161774820473339,0.0315788609121725,0.0177935894698342,0.0235128102329494,0.00656341341061273,0.0181538172126421,0.00289974871672105,-0.0064080946512004,-0.0270532163348416
"521",0.0338338804177445,0.0373935197791677,0.0181404553634692,0.0506995152601535,-0.0249866816607018,-0.00641783971868837,0.0796185049878626,0.0177616305798252,-0.0108621750688677,0.0238332003545942
"522",-0.0324975638123692,-0.0456816415591759,-0.0378617241585661,-0.0507488314161263,-0.0229970216368913,-0.0130218122123468,-0.0783031413611381,-0.0300324282445924,0.0237932057605399,-0.0121241352363949
"523",-0.0203431477166659,-0.00710561866527293,-0.0243055746928725,-0.00744974635553408,-0.00317138734987654,-0.000422361851259878,-0.0318193435249162,-0.0121341128517161,0.020223441340782,-0.00589103658931234
"524",-0.00301823452399053,-0.0128056964867851,0,-0.010154715371295,0.0186049384330653,0.00811090142208704,0.00638142077780879,-0.00465935877560486,-0.0270507288807519,-0.0192592500730235
"525",0.014046753770792,0.0335748902474333,0.0189798356228796,0.0298842192811086,-0.0238160106062602,-0.00861284649584793,-0.00380452357279304,0.0144684768567789,-0.00416473454141086,-0.0115811681446749
"526",-0.004896216842741,-0.00996690268850675,0.00931312056185174,0.00736252454992603,-0.0034991653440144,-0.00508574802444473,-0.0235517710325422,-0.0151009712618817,0.00802530792330391,0.00560380148302553
"527",0.0148808438994663,0.01938855479686,-0.00346015588969195,0.0210661901780422,0.000878050995957835,0.00234288315792908,-0.0153195264500338,0.000426136260400556,0.0105405135680645,0.0222897741548633
"528",0.0284969168436255,0.0263349762798082,0.00578695023275122,0.0501050912892143,-0.00311799618565878,-0.006056477098348,0.0685202713867143,0.0400166604243888,-0.00588112497066828,0.00743300010297254
"529",0.00137955321273675,0.00819678256566636,-0.0184120400176451,-0.005212339881002,0.00322522317086182,-0.00203030488402678,0.0136310422885546,0.012280439775505,-0.0141756452361044,-0.00541064938474589
"530",-0.0458092859907758,-0.0516083240421388,-0.0351699610209232,-0.0604595921471269,0.0217309774759527,0.0133881067260713,-0.0858803334152376,-0.0477155736678019,0.0213994451992754,-0.0128586343260043
"531",0.00589600242265265,0.00782711712856354,0.00486041477770871,0.0300299846055105,0.012971009203061,0.00771557085774366,0.0254099307704541,0.00127396463300911,0.0230573331455197,-0.00601204533501087
"532",0.000717611221212167,-0.00517776236577461,-0.00120935390639276,-0.00624727035139583,-0.00941577816521189,-0.000313639030577018,-0.0146727702543481,-0.0029686143692097,0.00953512829629299,0.00151228372584122
"533",-0.0107576666701107,-0.0115239349503811,-0.0266344248856129,0.00502916058487624,-0.0266131746929767,-0.00786925408816985,-0.0598942160861526,-0.0110587895803168,-0.00665444899977352,-0.018117878429032
"534",-0.0427742845526574,-0.0590451345558001,-0.0335821171075715,-0.0638032281230563,0.0311492545771381,0.0168150486012215,-0.0630062097426057,-0.0692477051381304,0.03133434798484,-0.0558688131967552
"535",-0.00239837347553906,-0.00439617715157814,0.00772204875753979,-0.00712681274627536,-0.00852311135136474,-0.00728006010333138,0.00413253558762716,-0.0189467277820532,0.0152960402921751,-0.00597174427432889
"536",-0.0107553888973579,0,-0.0140484770670707,-0.00942134814970297,-0.0170007711069867,-0.00555341609007942,-0.0385333020784626,-0.0254350631064896,-0.0117635636461226,0.0245768480119914
"537",-0.00972140543456845,-0.0124446664979653,-0.0129534484847275,-0.0253622369611066,0.00971666381440195,0.00284572956171902,0.0642022135552041,0,0.0211966802087298,-0.0111942597399849
"538",-0.0357785642603852,-0.0402439664259051,-0.0419945645200615,-0.0246282895094856,0.00923762319731236,0.000944454683690532,-0.0760512993008026,-0.0362497159070082,-0.0007157463993126,-0.00970331719433548
"539",0.0379099366351885,0.0427781993499088,0.0410957699450722,0.0547883000143483,-0.00104832160093582,-0.00377854038833048,0.0823111707860522,0.0275828171062134,-0.0306968168209306,0.0190527660614423
"540",-0.00787306604537819,-0.0288382182470822,-0.0263155964081334,-0.0171638462423863,-0.0115497892392524,-0.00905987008293363,-0.0252282361038576,-0.0278184197066988,-0.0166789923990607,0.0117521957846016
"541",-0.0162610156604223,-0.000836357876551896,-0.0121623454404237,-0.00873153105659408,-0.0105250238250261,-0.00255100096332772,-0.0423858476770782,0.0115462678349969,-0.000966226495625944,0.0211193055324381
"542",-0.022348889216779,-0.00711600084856334,0.00820785339947161,-0.0157629942861351,-0.00575725721192288,-0.000852821633351653,-0.0152761170825703,0.0143918551043265,-0.0046206856785016,-0.0118925004637856
"543",-0.0450425303116158,-0.0619731228792535,-0.035278000481326,-0.060762772691306,0.0165547241614432,0.010032215500227,-0.0700081555865262,-0.0631115802073938,-0.0183525537629025,-0.0502355994577631
"544",-0.0075070487444463,-0.00898864112431474,-0.0028130245993514,0.0140424636839713,-0.00668092397160824,-0.00127038717820116,0.00384957842216416,0.00574421922035651,-0.0097877378203014,0.00661170746738571
"545",0.023690701416953,0.0380955863010026,0.0267984613841856,0.0702273714345754,-0.00458128053664497,-0.00508923271725714,0.0264170579408491,0.0150569014703477,-0.0116615169739948,0.0350300751350248
"546",-0.0408475916710994,-0.0397556965685124,-0.0192309770261865,-0.0411274576786028,0.0278106213199945,0.0117233200390312,-0.0643422032891465,-0.0424550160522906,0.033711653752369,-0.00846112494133433
"547",0.00174409175756995,-0.00136495182735297,-0.00280120558086638,0.016867409864932,-0.0066695444781919,-0.00474060675233279,-0.0146407232185853,-0.018696359685435,0.00326125672923716,0.0240000562089202
"548",-0.0117526813184653,-0.0241456454873755,-0.0351121809551691,-0.0194313322858085,-0.00585055841891124,0.000423516371648391,0.0211615634727242,-0.0446383543121378,-0.0186369160403412,-0.00572919525600046
"549",0.0596093583072805,0.0732959327493279,0.0509463040189015,0.0811986745514368,-0.0191985451273721,-0.00729990725573082,0.132275393976095,0.0717947017019889,-0.0268300872253504,-0.00261919038814651
"550",0.00651268639913494,0.00521982290269563,0.00415489506231936,0,0.010820263095251,0.00714025934369178,-0.0171342186433115,0.0159494560754148,0.012253256322365,-0.0315125524628562
"551",0.0393718668083127,0.0359149597885933,-0.00137924830343894,0.0384442685652664,0.00476774910289746,0.00285676566984816,0.0788428538532784,0.0387228378153928,0.0210714747694298,0.0466376618266351
"552",0.00781482442298786,0.00167056041925284,0.0096684890829446,0.00559635717045071,-0.00503682958060048,-0.000737947949652873,-0.0212998701749726,0.0292195005415563,0.00219544461460908,-0.00880838321565069
"553",-0.00302297555781617,0.0104254357708073,0.0177840877934181,0.000855888896499346,-0.0157683405151126,-0.00570248707101451,-0.0735456332187249,0.0234947393430689,-0.00547645107963468,0.0219551233768189
"554",0.0305829957719235,0.0222868277115527,0.0349457490291181,0.021813499012489,-0.00544002397058918,-0.00191208769085716,0.0745238644391557,0.032520199137718,-0.00837006580275113,0.0214833462568833
"555",0.0223842396757592,0.0270485898557749,0.0233767900084092,0.0209290845157286,0.0378874898431374,0.0342626282327925,0.051639931451376,0.0310332069066936,0.0338737779445382,0.0125188655265474
"556",-0.01238630886244,0.00353787403199135,-0.00507625823379754,-0.00655983664184301,0.00124637745286549,-0.00339510264780785,-0.0569897327283686,-0.00628989639554345,0.0135353104967368,0.0207713816451687
"557",-0.02129379197618,-0.0117508022114509,-0.0216835088128814,-0.0136194874419436,-0.00555054627023877,0,-0.0744962409243519,-0.0134089416030865,-0.0080551353058852,0.0135659568000472
"558",0.0718292492698618,0.0729292522806639,0.0782270319734968,0.092468793243595,-0.00866113215107167,-0.00340686886411434,0.149897706044111,0.0411023221699049,-0.0161341389522017,0.021032562538039
"559",-0.0197033879252028,-0.0369414759412409,-0.0278115683462257,-0.0310228305876433,0.00951300005735645,-0.00144965375454509,-0.0714284661892787,0.00897265566973826,-0.0122719914797569,-0.0163857844833152
"560",0.0105460097006405,0.0149595626538377,0.0298508665609725,0.0150199157324626,-0.013461401329282,-0.00601619016803723,0.0138824523063985,-0.00222385677988468,0.0113249701371623,-0.0152308792253397
"561",0.0203809439686902,0.0120939783276619,0.0108695122001823,0.0272586238038977,0.0115980341858954,0.00260851262879536,0.0248256078827713,0.0160430294353899,-0.000543629032062398,0.0173997215694346
"562",-0.0180485888954615,-0.0403287920662756,-0.016726407135786,-0.0295678496428257,0.00741895271410908,-0.000624148276913483,-0.0401209258475504,-0.00350896143993307,-0.0134885021211791,-0.0185273076455011
"563",-0.0345548305573905,-0.0412452800397642,-0.0388822562121424,-0.0515623728179635,0.00382581590013942,0.00427029865935746,-0.0548110219112045,-0.0528165710296815,-0.0078288563716209,-0.0363020355662409
"564",0.00926488582588814,0.0381494699001119,-0.00126416575881039,0.0218285353234036,0.00714576084321505,0.00176270659467126,0.0621610595540842,0.0250927538020804,0.00333402967323759,0.00452038323437498
"565",0.0193665046949976,0.0234558353865921,0.0291138364487624,0.0330511267288476,0.00912582345189294,0.00245043460394267,-0.00903384528820761,0.0117857262415813,0.00830748790770364,-0.00249996577856626
"566",0.0292377743177543,0.0469824580487674,0.0356706843733832,0.0542333358298159,-0.0122213093479184,-0.0065249915099338,0.0661914053815125,0.0640685085140178,-0.024497374761039,0.0385963742912467
"567",0.00994815642990976,0.00839116103193915,-0.00831366477124462,0.0122130868897814,-0.0204625885742407,-0.0114674186941283,0.0895906929308636,0.00505255173874386,-0.0136262044946103,0.015444053609444
"568",-0.00783262264018791,-0.0188132488306051,-0.021556961918403,-0.0124313566208982,-0.00427486968864377,-0.00232067116950818,-0.0160353103264843,-0.0146624286546015,-0.0264870316925234,-0.0123573436304513
"569",-0.0233256561761981,-0.0265487114022118,-0.00612008162273048,-0.022954571931514,0.00253708778813611,0.0025370567268832,-0.0752428256634814,-0.0153062721533518,0.0172393696694981,-0.0178056351805647
"570",0.0107779810668835,0.0102271337996247,0.00738946224119719,0.0147784213545288,0.00885711172124348,0.00495558368974947,0.020997227505805,0.0250428197890273,-0.00149869729072394,0.00734928855250017
"571",0.0397425110781291,0.0217475518956474,0.0366747087938986,0.0436893155428499,-0.0125425438695808,-0.00587593964181943,0.119353840542958,0.0421230491946196,-0.00346383785401416,0.0145914913061271
"572",0.000233522907074013,0.0176144951543995,0.00235834881960484,0.00608222376276757,0.00918513837751478,0.00591067038423998,0.0127949452309573,0.00525496110358836,0.0181902333029831,0.00431451718146958
"573",-0.0172437182292511,-0.00937619688194513,-0.00941148404723169,-0.0160027920689488,0.005227788775239,0.00514117155047877,-0.0819562196502126,0.0072375579322892,-0.00580330015259334,-0.0181385200973956
"574",0.0106698761951873,0.0152896249157992,0.00475062978892105,0.0144561790904019,-0.00173401218682279,0.000939664070061408,0.0818631399949221,0.00518992843483002,0.00148789052920151,-0.00631979731497179
"575",0.0146628837743603,0.00609521607175711,0.00354568959863255,0.00855011466602296,-0.00791084663484753,-0.00396315578423034,0.0407695624624218,-0.00198576323009214,-0.0193143085714287,-0.00440312116309871
"576",0.00670550218936583,-0.00178190925340571,0.00471160462720799,-0.00706479654560388,-0.010989129774283,-0.00806155542147236,0.0100281477876529,0.000795663666328439,-0.00687562071729675,-0.0073710074952722
"577",-0.0419154194157503,-0.0485541984014617,-0.0222742073584838,-0.0487370767670942,0.0151427084960614,0.00696621942319386,-0.107043014485229,-0.0588467973834165,0.0203003517918288,-0.0376237562217255
"578",0.0195373087832136,0.0228894266688719,0.0119902282837701,0.0213163079095244,-0.00988011426447277,-0.00387863246657261,0.0913827032731684,0.0190115150145342,-0.000690028775964135,0.00360077366973188
"579",-0.00611340278583294,-0.011005062171634,0.00355487833837853,-0.00842165580888243,-0.00606524849414614,-0.00241999081744004,-0.0337470587276314,-0.00373153378570878,0.00563929112256067,0.00153775748535745
"580",0.00981788317619503,0.0315280031082243,0.00590295590451984,0.0155094062166232,-0.0000986411377825736,-0.000211372009990884,0.0415155617274297,0.022888214574041,0.0162509275435201,0.0133059086425964
"581",0.01511037202069,0.0172601603951548,0.0152583065577649,0.0189092139162104,-0.0100401630378709,-0.00390350235069647,0.0528310344995166,-0.00325508033037558,0.0103603374878263,0.0151515687072972
"582",-0.00946220729432889,-0.0130788232184269,-0.00231245243510991,-0.0335473972232342,0.00427542529258251,0.0041310445905296,-0.056490261829504,-0.0191834296398533,-0.00791349745972469,-0.0248755890277783
"583",-0.00314513962402685,-0.0028653507420916,-0.016222520594297,-0.00332380344533134,-0.0163364567887706,-0.00485275642987582,0.0108280720311185,-0.00457782870016898,-0.0141557349925686,-0.00714296929139702
"584",0.0212691109875147,0.0312499777346054,0.0082454412208659,0.0526123367603448,-0.00885791229982902,-0.00540572581009646,0.0396976624898386,0.029264182055893,0.00660970940170924,0.0231244135623185
"585",0.000343170055334241,0.00452802340302094,-0.00584131494036633,0.00915158637234725,-0.00396027738576787,-0.0017060526744056,0,0.0125917017093071,-0.0120005091814669,0.00351577321474195
"586",0.00537609137652151,0.0124827070535571,0.0152762366857619,0.014649500031656,-0.00688285736075189,-0.00321104830989949,-0.0339393933124374,-0.000401284618166686,-0.0036667813796305,0.0300301367672682
"587",0.0340199161562,0.0410956617593292,0.0266204943188155,0.0690959857665323,0.00329540842752585,0.0009655919071625,0.0865744777276747,0.0389247823754435,0.0194364814066641,0.0194363296856011
"588",-0.00341085918194717,-0.0108550664900087,-0.00338247579409712,-0.0090032667078499,-0.00123140200980421,-0.000213769625158733,-0.033486949178387,0.0023174958543013,-0.0043998082626332,-0.014299382269237
"589",0.017334444857247,0.0216163897250787,0.023755815201091,0.0171967332435083,-0.00236360490833976,0.000429107156572295,0.0334526150021266,0.0354525119361275,0.0146175750708215,0.0265957801542649
"590",-0.0138918242786343,-0.0179037301786209,-0.0232045716843375,-0.0248804593188136,-0.0244126392395587,-0.00836873842028663,-0.0578037067024944,-0.00744340481339112,-0.00111680811797177,0.00188410047824861
"591",0.0233327739755311,0.0477293210159619,0.0407239234315506,0.0333661408019605,0.00242838800074074,0.00118971911762733,0.0677919696998113,0.0292470386261785,0.00603757812974992,0.024917674809716
"592",-0.0187138944497452,-0.0306863654865186,-0.00978233312086352,-0.0234252145387934,0.0142192056326029,0.00940291270896565,-0.0293017702587298,-0.0280512397305789,-0.0032229494368875,-0.0082568156770203
"593",-0.00295952217094764,0.00979114936770853,0.00548816000146091,0.00713142130568434,0.00363496990313572,-0.000642550348881277,-0.0159813940971858,0,0.0112609541473752,0.0101757669694855
"594",-0.0251730874411751,-0.0303814713272572,-0.0185588100082349,-0.0366915406069922,0.0108647388808747,0.00460628213268022,-0.0679699658519586,-0.0431034368559238,0.00429987886328154,-0.0114468713857856
"595",0.00857063057273577,0.0103335053852536,0.00111226344454352,0.0143670209856757,0.00389045265899024,0.000106369914119275,0.0319456940075982,0.00940033560396691,-0.000658656302937932,0.00648449018123598
"596",-0.0081617315190895,-0.0131972485304644,0.0100003543018643,-0.0092227550835714,-0.000305844884208817,-0.00245203249723391,-0.0328326966909558,-0.00388045641813184,0.00571244650897995,-0.0253106155559778
"597",0.0284069762870887,0.0434636770257879,0.00880101198375294,0.055518598338584,-0.0155046022001931,-0.0058789565357148,0.0750078689546387,0.0268796567362333,-0.0129983829711071,0.0264399184207804
"598",-0.00120563173455601,0.0124962269352764,-0.00654330391688474,0.0113384242175043,-0.00528391268744899,-0.00139880493104316,-0.0159396572950115,0.0170717748593929,0.00664008403452754,0
"599",-0.00669431791738229,0.00474691561008034,0.0131720074726422,0.00311464139127637,0.0105201246001814,0.00312363413158656,-0.0116138788161406,0.0104435564417544,0.0141820691972523,0.0160994686754468
"600",-0.0143634894829265,-0.00440965978601904,-0.0130007613470291,-0.0186278866970494,-0.0251495635159146,-0.010948172957299,0.00185539100989662,-0.0103356158542205,0.0173441517615176,-0.00814846504239086
"601",-0.00212990616936604,0.00379638540613492,0.00329296878463436,0.00442892274245366,-0.0111017179632918,-0.00586172374186533,-0.0212965954470137,0.00522132722720281,0.00319663299300221,0.0146050497443448
"602",0.0256119515928412,0.0211157762178269,0.0328223657416218,0.0119685037223443,-0.0150749524999133,-0.00665938479919548,0.0517186260348024,0.0330241735984416,-0.00414232598741737,0.00224927486095283
"603",-0.0178528008239875,-0.0169753896229066,-0.0190674232263711,-0.0115157578539681,-0.017694232295954,-0.0113201827162321,-0.0332828734363888,-0.0114940063430413,-0.00330636725029088,0.0044882691767838
"604",0.0139400198061812,0.0128726256822698,-0.00647964522313393,0.0308563205282217,0.0144762385787418,0.00522535380551958,0.0189205471495413,0.0148987119971011,0.00845372953837553,0.0183200938637791
"605",0.0177080807996977,0.0136393297991024,0.0184785120168689,0.0152722171197459,0.0258165278548323,0.0112784728525641,0.0273968461463647,0.0329390201545616,0.0207979524787341,0.0193066290542936
"606",0.024208299143319,0.0284405368282232,0.0160082652523275,0.0421177020046155,-0.0295628252894674,-0.016318741988639,0.0420742989858205,0.0183708017487589,-0.00488559266794986,0.027550648242207
"607",0.000843737119398336,0.0071363690750037,0.00105056296485673,-0.0144342415812048,0.00537869723226825,0.00334392615064982,-0.0147852998526596,0.0139551834302751,0.00658098798973183,0.00418930158616559
"608",-0.0126513706622108,-0.0345438921663627,-0.0220356964557118,-0.0354419923914093,0.00939156032213884,0.00611182528232179,-0.002308542866999,-0.0184624493603156,-0.0202365813591056,-0.0333750258162775
"609",0.00939662844930944,0.00795104327925489,0.00751097360668762,0.0185237655712804,-0.0206625529383349,-0.0115963176932051,0.0295051029570907,0.00273523445752866,0.0192776074874437,0.0366854001460537
"610",0.000211473219034808,-0.0127426853457765,-0.011714798055897,0.00208712931859933,-0.00762217504292817,-0.0099459239625912,-0.0126439425661554,-0.0225097925762945,-0.0261873004410069,-0.00541225372086029
"611",-0.00412447342724931,-0.00522433485902984,0.00538798062562718,-0.0154715342736115,-0.00255936139500512,-0.00507843297969757,-0.003699833488505,-0.000348864182597941,-0.00160069364636317,-0.00251151998290522
"612",0.00509746077336515,0.0120481516376085,0.00857452416247728,0.00181338436147183,-0.000112081928305918,0.0043099833988034,0.00114302313552583,0.0150087973672113,0.00288589146827478,0.00965169779847508
"613",-0.00253590438887197,0.00274718692297515,0.0010626512980132,0.0126696001018634,-0.0157367628315676,-0.00598596043431998,-0.0191158207936847,0.00447081925594373,0.000319716501764544,-0.00374059749461575
"614",0.00444963739222293,0.0167430266538091,0.0169849162144335,0.0214477609274719,0.0111129781805264,0.00681773378925588,-0.0186155948648185,0.00581946390396992,-0.00170470912311205,0.00917814283389506
"615",0.00274171551190139,-0.00508990013255117,-0.00104344844184301,-0.0160397171048318,0.00897068772183451,0.0053053472582647,0.0281564936745675,0.00646686635596616,-0.0163286984950489,-0.0140553730163712
"616",-0.0229280195871653,-0.0373156569834173,-0.0177641751905652,-0.0358624678306821,0.0090039635606276,0.00449063562467722,-0.0449695174114619,-0.0246868745023227,-0.0116089836521425,-0.0192872499722414
"617",-0.0135630856673975,-0.0128164670841014,-0.010638365067936,-0.0150630451435095,0.0174039041273997,0.00558852586310188,-0.0141866642835893,-0.0149099153110465,0.00911088933284065,-0.00384783372232922
"618",-0.000982095558690999,0.00316636008793569,0.0118282366706417,-0.0112359166666336,-0.00562968657533292,-0.00266750306333563,-0.0140840419674385,0.00457599349010462,0.00456867181551179,0.00300442766130105
"619",0.00731825109765483,-0.00315636589693669,-0.00850162675841681,-0.00284089927416109,-0.0151349700467472,-0.0121476763830832,0.00496857653877147,-0.00455514915721467,-0.00801296173281996,0.00128359132876055
"620",0.00368597362150114,0.0145659742473865,0.0160770591737365,0.0050647958129022,0.0137087056075984,0.00462559562857945,0.010815649266706,0.00997142033827703,0.00316560415712686,-0.0085468920092806
"621",-0.0299871089995931,-0.0362212911920808,-0.0221520467293371,-0.0362205108278578,0.00970728245456498,0.00538956182469019,-0.0510546268971652,-0.0278561352190982,-0.0147987047921936,-0.033620804004005
"622",0.000783938047397958,0.020198613736957,0.00650780292277764,0.00649004302928868,0.0117732923011045,0.00324013192271422,0.00869856381688794,0.00652895382691088,0.00419700680144675,0.017395175235059
"623",0.0086184907866278,0.00194735411203673,0.00215498333395137,0.0219314725074216,-0.0100350140247463,-0.00378576554495302,0.0164380391175385,0.00504490016803527,0.00582928961349061,-0.000438398234711701
"624",0.0217479715133455,0.0129576223879935,0.0236561315674853,0.0297887264788514,0.0183321023225167,0.0125168932688606,0.0159492281830158,0.0340627048943116,0.00940405717017123,0.0087719456635289
"625",-0.00260593609031756,-0.00319780136754266,0.00315103119118154,0.00528766478346454,0.00169496017339776,0.00132431427023194,0.0087909455161701,0.00970826623312826,-0.000216628755641324,-0.00826089106396555
"626",0.00936387032400932,0.0112286549241993,-0.00523544202653214,0.00742594061497748,0.00147940811324743,0.0020941060079287,0.00248967499921848,0.0058380889688241,-0.00270885250071673,0.00964489652745826
"627",-0.00809063120923637,-0.00444178233121251,-0.00736826401212143,-0.0101353452735408,-0.00168836514521842,-0.00263990813106185,0.00651952219119045,-0.019119171660954,-0.00934377434437439,-0.0178027572355389
"628",0.00413269303758002,0.0152965161342971,0.011664685132146,0.0183057943707314,-0.00198369000473553,-0.000640619210295457,0.00987094259778787,0.015662969882217,0.0132704430796227,-0.00397881616864659
"629",-0.0272929980810944,-0.0310735514956501,-0.0220125191320378,-0.0274221154767249,0.00233818799581753,0.00331929816600574,-0.0455103251470516,-0.0215895785511684,-0.0123389870368978,-0.0221926019969989
"630",-0.000111578102719556,-0.00161952886074035,0.00643113956072461,-0.00219283646260304,-0.00190897533864898,0.000662142708579783,0.0208001826656714,0.00910628971919047,-0.00536984109589045,-0.0299592023076115
"631",-0.0193767696263193,-0.0295263412415536,-0.0106497758671972,-0.0235481275111185,0.00669414875557761,0.00396835359557879,-0.0369905445091565,-0.035751203876707,-0.000550936523778467,-0.0159100812892855
"632",-0.000681003458896434,-0.00668677944815999,0,-0.0115756284950791,0.0184688350249707,0.0115281718231601,-0.00976574677157505,-0.0104391386127212,-0.0158747879602555,-0.0123634141565601
"633",0.00193172924666452,0.0151465352993103,0,0.0178921002844827,-0.0119164241076553,-0.00586149286857818,-0.0161076480940402,0.0080029566911759,0.00268852927148622,0.00625904125719567
"634",-0.00238184927957796,-0.00795784229121255,-0.0107644467361558,-0.0118248906242308,0.0092287001861906,0.00622333656668128,-0.00167085777065823,0.00360872979664673,0.000782035509282908,-0.00765554569948457
"635",0.0243290308740756,0.0257354744295135,0.00217647928014575,0.0071151762208721,-0.00561218188356871,-0.00358068728553873,0.0394913535880483,0.00898968173589965,0.00680955555236551,0.00530393685595221
"636",0.00566099774098272,0.00260675999440863,0,0.0109185349673826,-0.0166146534877774,-0.00664243989651159,0.0115904297174223,0.0242335246641401,0.00687433181340857,0
"637",0.0292461069655889,0.0425738290768329,0.0108577535470193,0.053684815455401,-0.025717522004662,-0.0129359809610767,0.03437318445495,0.0208767133348,0.0157471647560217,0.0263786816745606
"638",-0.00160852261601263,0.0109102249505535,-0.00429672207108922,0.00180891161806529,0.0107976453732268,0.00599745095452353,0.0129233046496309,0.0248805901368225,-0.00281867959277282,0.00233656119252856
"639",0.0109546716809117,-0.00370019589900761,0,0.0102317750875882,-0.0154307258168292,-0.00673432994498624,-0.0233903118055084,-0.00897866281286563,-0.000543629032062398,0.014918402839005
"640",0.0106235598444955,0.019498357807082,0.0129454026319791,0.0357463606488122,0.00525998262303817,0.00366815800078224,0.0323483049770039,0.0218116551800343,0.0146850756010006,0.0165364813130622
"641",0.0046253467176891,0.00455398140312124,0.00851978238509665,-0.00287634842904239,0.0199525040881154,0.0111846651846708,-0.00210909873345388,-0.00426880186260048,-0.00160808320763384,-0.00361499950632049
"642",-0.000208904442373647,0.00392856794391561,0.0116152861537862,-0.00230744704232588,-0.00897889826831133,-0.00591413146066044,0.000906067035391755,-0.0042879515976233,0.00332873413493195,0.00544224272584604
"643",0.0220825315106481,0.0174596098159265,0.00417543720213165,0.0283315360549901,-0.0183367110568834,-0.00969516054162456,0.034690568773236,0.021530442234643,-0.00192636982178152,0.0207486147016711
"644",0.00409588056676857,0.00739622004136908,0.00519715802525078,-0.00477905293023329,0.00483457806225807,0.00211408103492916,0.00874619873387839,0.000648506884140865,0.00160842801611771,0.000883861571832734
"645",0.00295727849015925,0.0014683997986733,-0.0020680094918073,0.00875704078662776,-0.0114815068732073,-0.00466241564147529,0.0187864262018251,-0.0116657374526016,0.00321159391021975,0.00397354664689109
"646",-0.00467758744406654,-0.005864865142723,-0.00103628729574223,-0.0044803158231419,0.00884986277717204,0.00200747090569187,-0.00397164322450838,0.00557387862200387,-0.0170739303924227,-0.0109938289580486
"647",-0.00245156275843261,-0.00973465427540232,0.00726144281983432,-0.0225034269570237,0.00548206491323544,0.000667859026830087,-0.014241149528304,-0.0091296608952266,-0.00987953523092455,-0.0257892071251772
"648",0.0104454523610242,0.0196603271626243,0.0113288150574948,0.0247478994054577,0.0141770441792075,0.00400455081915596,0.0349609902572365,0.0164528061807874,0.00460532909885947,0.0310360066831867
"649",0.00141885907242667,0.0169443202013173,0.00509152227489484,0.00477382532804449,0.0194617787587175,0.0100812960882311,0.000837557178522852,0.0213665087663568,0.018882284908897,0.0199203653748934
"650",0.0164966102170938,0.0264292518081037,0.0172235062895134,0.0374510257486564,-0.015154262768724,-0.0106258407830579,0.0198048023278308,0.0288430339051875,0.00557048753230815,0.0282116866853799
"651",0.00258818363586677,-0.0033586803397655,-0.000995913904622281,-0.00915933256883672,-0.00795230252792289,-0.00289098321570436,0.0475930039872501,0.00462117411591945,0.0086289227028149,0.00042220018779604
"652",-0.00287946340479417,0.000842412219705047,-0.00697861614724127,-0.0084284734084682,-0.0149476963789874,-0.00568696226118581,0.0404697786622834,0.00275993898275106,0.0010561787072243,0.010548596042903
"653",-0.00517866511040266,-0.0084175759003462,-0.00100412333739364,-0.00822577839172611,0.00340894595145014,0,-0.00627336300005044,0.00152882313173341,-0.00189914540936009,-0.0229646233327346
"654",0.0131140119903752,0.000283171655858228,-0.00402001829622767,0.00995284551704634,-0.00832906693011992,-0.00661644742519452,0.0464647105645717,0.000915916095461045,-0.0089851798939784,-0.004700702637916
"655",-0.00207490144718026,-0.00735489101310738,0,-0.0112236812384523,0.0124879727830669,0.00643462131074624,-0.0197878220275276,-0.00274551432317161,-0.00874666666666657,-0.000429451290466343
"656",-0.0124762893080759,-0.0108293247136905,0,-0.0188263129465797,0.0115690130528179,0.00695483029203969,-0.0295418718138504,-0.017130468997643,-0.00150649951576454,-0.0150343792638081
"657",0.0107290987629125,0.014693094638345,0.00504543364630727,0.00902975504691872,-0.0106822225770986,-0.00278424842342673,0.00659550726097136,0.0289448400765642,0.00172428061510632,0.00523324715238638
"658",0.00763836615574487,0.0167518905378488,0.00903617703221449,0.0173375500198363,0.0141786283164393,0.00781910260408281,0.00478861607812697,0.00574694585403557,0.00828406696990003,0.013449063960312
"659",-0.00767939541902418,-0.00949469838420303,0.00397986842184528,-0.0181414895063631,0.00387129028951305,0.003104124096595,-0.0090298477592673,0.00330842924536001,-0.00768246897479219,-0.0282533912361369
"660",-0.0246055895669929,-0.0352410165472904,-0.0277500987532139,-0.0391939056249633,0.014783223676845,0.00684979501592009,-0.0501138266527033,-0.0344723403676045,-0.0149462258064517,-0.0149779951796416
"661",0.00793425136747028,0.0187024507187368,0.00815483777916404,0.0218531954777126,-0.00580596625477992,-0.00351129146791962,0.0122573787650881,0.0229741181348635,0.00491209469586185,0.0196779575566206
"662",0.00877987171471295,0.00975328930893316,0.00303314601083149,0.00256613019214269,0.00828236210581457,0.00374414835586778,-0.00737074331496146,-0.0145676040132027,0.0051053770390046,0.00701749333334312
"663",0.010304111813515,0.0090909187533581,0.0120965904468884,0.0173493595851926,0.00821367641709125,0.00263315930469066,0.0405728025206897,0.0163224960056281,-0.00280992113703582,-0.00827519375240693
"664",0.0196057877186682,0.0295606956562038,0.0109565458065608,0.0150966401633679,-0.0205765192550476,-0.0101773456990831,0.0221712767247502,0.0148488450663045,0.0149561617521241,0.00746599767470402
"665",-0.0000970250465600619,-0.00136698673791347,-0.00197021124240437,0.00440621052750179,0.0181295797753116,0.00619161885109087,-0.00573414817573936,0.0050760752498975,-0.0139883179073504,0.00174365530253318
"666",0.00194237381033924,0.00766684903181858,0.00789690561182432,-0.00219331932907663,0.00565580061147331,0.0026374383097989,0.0110332809103484,0.00950702971359174,0.00454847323146956,-0.0143603410888363
"667",0.0000974189722937613,-0.0040758560700358,0.000979771826582043,-0.00302317190307833,0.00458283010415883,0.00131478937490415,0.00446402236810717,0.00176574016079001,0.000323404477718725,-0.00264897051125457
"668",0.00222924695599014,0.00818548920983586,0.00293520652800772,-0.00192927490829287,-0.00393973097982947,-0.00273656606443295,0.00790136184877421,0.00793193320529606,0.00431082008502193,0.00841077740029217
"669",-0.000193814338504961,-0.000812124353579025,-0.000975948203825183,-0.00524716406123438,0.00458041115030094,0.00230507481220243,0.00661461456813428,-0.000583240453737921,0.00729693084457694,-0.00219496822668053
"670",-0.00889915822437248,-0.0062296083753427,-0.00195257371170676,-0.0197113827591793,0.00093195299743587,0.00295589499904092,-0.0124120503713809,-0.00670747979142272,-0.0050069349630254,-0.0272766279455596
"671",-0.0220574510120475,-0.0283454768952062,-0.0146774992020436,-0.0189746893647958,-0.00241953768136549,0.00259478193680818,-0.051010402279012,-0.0284788199646797,0.0053533189431838,-0.0153776794646028
"672",-0.00379252677314201,-0.00364669350415825,0.00297940605788649,0.0106815359002139,0.0145745116064186,0.00546006936674814,-0.0197351786604115,0.00604388405672762,0.0243876459129362,0.00229675452761691
"673",0.00831517976231289,0.00760146663775174,-0.00297055556663606,0.0199939627312258,-0.00615656775619777,-0.00358444111414913,0.0177482475976809,0.0156203245314357,0.0132030041957998,-0.00504131910971206
"674",0.0140092433184216,0.0192791173114086,-0.00198562572840821,0.0193225000723072,-0.0170345248405753,-0.00599419721319516,0.0119731973781436,0.020112127142611,0.000718243389270068,-0.0041454986395717
"675",0.0086217070039265,0.0249451516463586,0.00895513644628276,0.0206043712086315,-0.00703733627953163,-0.00230201117426954,0.0321499910145258,0.0171067443297406,-0.00102531529811656,0.0185013728514223
"676",0.00767472375140832,0.0117679008747673,0.00394478098894502,0.00538367806337936,-0.00116383668043374,0.000878366179964729,0.0201843977552796,0.0188141451763855,-0.00359230216565753,0.00408723115819432
"677",0.0102190556655668,0.0113666049593897,0.0117877247238389,0.0131189108374088,0.0184260977400899,0.00746665625462128,0.0141670394756346,0.012590749108212,0.00638643373740355,0.00542728758512201
"678",-0.000191159527903273,-0.00313636549495988,-0.000970977654562999,0.000528477506621883,0.00551164332657272,0.00294362586025954,-0.00313125492589217,-0.004420897483848,0.0110542685072959,-0.0130453034291789
"679",0.00486799031341967,0.00498175090991126,-0.0038872776299812,-0.00369738855966617,-0.00992722751981234,-0.00586849498329434,0.0287513942829145,0.00471832954478302,-0.00830127564589267,-0.00546948107058731
"680",0.00417941837547819,0.00391319705697901,-0.0078048950539098,0.0119298063093556,-0.00511846579980235,-0.00207716390005519,0.0176135846366765,0.00414333115109122,0.00959578409142292,0.0233729683713699
"681",0.0151342797973077,0.0184511883981964,0.0049166527075839,0.0251506484863799,0.00178527692393216,-0.000766826445377955,0.03900323356852,0.0198076366020228,0.0102123557085469,0.0129871590421937
"682",-0.00149070671331197,-0.000765563989810314,-0.00978510701590951,-0.00536688497992099,0.0125754990428066,0.00493283231706765,-0.00488661094676635,-0.012139265808443,-0.00570521446480976,0.000441898573175337
"683",0.000637031648793362,0.000766150527064635,0.00494085631892571,0.00282639130963025,-0.00890079846257541,-0.00534481491081584,-0.000223246638710206,0.00607254916678235,-0.00674449392971577,-0.00883775159514855
"684",-0.00252959067733904,-0.00918591929395562,-0.00983301066065201,-0.00871136121222116,0.00229703059528674,-0.000658227988538096,-0.015851968932063,-0.0148152447254841,-0.00314175540978534,-0.0218456740229847
"685",0.00582410691588575,0.0113311329916117,0.0129095887031254,0.0152495708139451,0.00208375372043035,0.0026342137946509,0.030923291617883,0.0158731710514459,0.0133183914872064,0.0164083024803074
"686",-0.00831196141839741,-0.00789410216496778,-0.0107840311323422,-0.0150205144157008,0.00301519139801854,0.0021887825011575,-0.0335256331144602,-0.0175438141604158,-0.00842777181554688,-0.022421542462665
"687",-0.0110190837971599,-0.020276937768582,0.000991097237334371,-0.0196435287750056,0.00290271326001368,0.00273041567384857,-0.0330806500922164,-0.0181360343415252,-0.0129515225548613,-0.0128440036923365
"688",-0.00533285955020346,-0.0044538088767605,-0.00792092748932238,0.00421858816575638,0.0127131819716666,0.00403019596849163,-0.000712765481475475,-0.000852737897565126,-0.00563816487017432,-0.00789966405563647
"689",0.0179035244131458,0.0142102298368736,0.0079841695171301,0.0128644407767267,0.00877704273371238,0.0017355299184898,0.0389919691672038,0.0145053468742784,0.000515494845360953,0.00889941747812428
"690",-0.00301000049802536,-0.00155655635501273,-0.0207920488229255,0.00233236949280613,-0.000910379008571716,-0.000432494241289216,-0.0167049828725467,-0.00616788418690983,0.00391547643744028,-0.00371406505878014
"691",-0.00386790957687777,0.00155898299990853,0.00505539490108609,0.00620685532075371,-0.000912041417540865,0.000757911818145551,-0.00698140358465582,-0.00310279932841606,0.0145745458277737,0.0279589470361863
"692",-0.0248132304880023,-0.0298388685708861,-0.025150525794192,-0.0272426640318921,0.0136966806365397,0.00752300919597371,-0.0424186375274697,-0.0200906580851326,-0.00971167445041321,-0.00634633504819593
"693",-0.00466119439349533,-0.00909340490127974,-0.0134160883424602,0.000264168949636989,-0.00692108207677433,-0.000430695760597621,-0.0097897093647008,0.00664169772813961,0.00490350398307782,-0.0100365005487431
"694",0.0149278875404701,0.0145748952119924,0.0083680302800595,0.023243862995656,0.000100985796375852,-0.000107979901912802,0.0269404740338377,0.00114785155615071,0.014740235394727,0.0322580997056205
"695",0.0143242663518754,0.0188882706204554,0.0114109542162824,0.0165204170939406,-0.00989705774326277,-0.00323435003937589,0.000240433182273181,0.015758791195704,0.0246443498296935,-0.0120535907304756
"696",0.00274855064591795,-0.0026113479708183,0.00923092702439354,-0.00101600603883611,0.0117304854299649,0.00638123837129645,-0.00312808796616426,0.0146686929189728,0.000782186163298615,0.00180756951475836
"697",0.0076562729553582,0.0172778515691752,0.0111787769601388,0.012201487410431,-0.0104854012455645,-0.00365416831631438,0.0188271290836857,0.00917448729638726,0.0125048650595461,0.0198466927695415
"698",0.00609689410904068,-0.00643332890699799,0,0.000753140744667036,-0.0229242777567046,-0.00959938881849298,0.00971342337632675,-0.00247938580543972,-0.00771905642337956,0.00398048486315061
"699",0.0039157235329057,0.00880563884746732,0.00200993383020043,0.00828148192178069,0.0015645808822784,0.00294058380394691,-0.00164220072670873,0.00386614076596326,0.00700118658114302,0.0202642210679891
"700",-0.00204314730276556,0.002310879683594,-0.00501519121690586,0.00174201246355166,0.00520503603810973,0.00228066117732473,-0.0150415708226476,-0.00687742745501507,0.00675940530628449,0.0112263661355538
"701",0.0172154426813984,0.0217724279753304,0.0110886293796415,0.0322978434068195,-0.0148112080593211,-0.00682620882798057,0.0367456113850961,0.0340719651153352,-0.000767331656103321,0.00768576514257147
"702",0.00365946804362371,0.00777123166909499,-0.00498492221894886,-0.00553528825270666,-0.00462559532184537,-0.00327249063784574,-0.00759511696305792,-0.00482190239171854,-0.0126703685928202,0.0101693954337263
"703",-0.00747414270434454,-0.0121888018741386,-0.0180362629580185,-0.0137948186688091,0.00813348789238311,0.00459642079919997,-0.0271338559006803,-0.01561220756091,0.00311101494156141,0.00251683053248986
"704",0.00826523219605768,0.0151094882462255,0.0163270599772483,0.0191410877033176,0.00785673148906429,0.00152555355009265,0.0231230905222297,0.0210555442424927,0.0101764198488079,0.0142258758004092
"705",-0.00528270151071308,-0.00297720669474644,-0.00301240010909509,-0.0132436345781558,0.00540620086735188,0.00228399681741487,-0.0186390467273391,0.00107083535436314,-0.00777132281191617,-0.00618816184932824
"706",-0.00897366578923575,-0.00273685614321462,-0.00302092851311431,-0.00536850368765729,-0.00599692528693663,-0.00227879206359416,-0.00783487073738376,-0.00642032914935131,0.00319089157205354,0.0211707498222049
"707",0.0101634070929015,0.00998029296896474,0.00201996394519832,0.00834165305447843,-0.00488893003865121,-0.00293695532134564,0.022493074948905,0.0123852822791561,0.00163853493975918,0.00812996973268176
"708",-0.0114332723384898,-0.0170455119210962,-0.0231850989533958,-0.00827264551574347,-0.00752603361107174,-0.00490891081792999,-0.0109990445093965,-0.0249995815358321,-0.00413779838602391,-0.00362906586020384
"709",-0.0108251097993148,-0.0160846669779047,-0.00309633688095767,-0.0125119065021637,-0.012954294162776,-0.00570242797414477,-0.00615211697884344,-0.0155487746788936,-0.0157502853560786,-0.0182111281800219
"710",-0.004583143806692,-0.00740707077313918,-0.00414067200319357,-0.017391337081498,0.0136580462518634,0.00860104920586369,-0.01523825567147,-0.0135768947183448,-0.0000982034154898281,-0.00700753571954482
"711",-0.0188875760827661,-0.0270202452779299,-0.0103950327451554,-0.0457649477498104,0.00473723055165487,0.00306114394355594,-0.0418281084598742,-0.0410112900929821,-0.010996514698017,-0.0257368123829955
"712",0.0214537575057294,0.0330600785992929,0.0157559746427494,0.0442502139183281,-0.01089592024389,-0.00479522108138564,0.0431490712502278,0.0330991434503654,0.0194579464074871,0.0311036398292528
"713",-0.02897336205054,-0.0358422211760152,-0.0124094209300626,-0.0466885640572684,0.0145109828760861,0.00744664517119609,-0.0191095888327565,-0.0221149154972435,-0.00155811663145167,-0.0252065640847321
"714",0.00733872292521243,0.00743480349015768,0.00942421626099565,0.0149053892220399,-0.00442010386974456,-0.0026307424132046,0.00147966952602596,0.0127573862562995,0.0138495856222527,0.0173801378940006
"715",0.003163575873391,-0.0076436646727529,-0.0010373312051235,0.0015733410793386,-0.00999498382137642,-0.00230803345076513,0.0142818663952748,-0.00314924948138284,0.0241462440831046,0.0141666878942486
"716",0.00257998391811642,0.0143424049049878,-0.00207672337222897,0.0185915932541181,-0.00913896575584905,-0.0027543956526801,-0.017965257001046,0.0103385067571848,0.00601163823043049,-0.000821681464220014
"717",0.0183950101269197,0.0172822683169469,0.00728386070039466,0.0205651779670062,0,0.000220863632895307,0.0207663991615701,0.00682203455995634,-0.00112040151485349,-0.00534540630864588
"718",0.00262037816958349,0.00205920409732174,-0.00619814492294046,-0.00125923054344423,0.000964861203544443,0.00298249976971854,-0.0154998114030002,-0.000564389758837103,0.00420636555786991,-0.0177759529768661
"719",0.022776069001921,0.0300539103705386,0.0114343023148926,0.0368221776626056,0.00117848346549709,0.000440399518840451,0.0469862418915117,0.0364406018918813,0.00707439262775766,0.0164141340305319
"720",0.000182467260581021,-0.00274306719156592,-0.00719415373072207,-0.0046218339376376,-0.00181903349913182,0.00077002097416301,-0.00493454419078287,-0.015262794232761,0.00184857192257004,-0.00496887633467813
"721",0.00511008023430803,0.00175053455060392,-0.00103518351660392,0.00855350864458071,0.00418151750307927,0.00286068329297917,0.018418098575504,0.0102403530961106,0.0111633823338257,0.00665829530987594
"722",-0.0101680184504956,-0.0107340033695977,-0.016580410349267,-0.0222923746287402,-0.00181521079369318,0.000328731736832788,-0.0118245543091517,-0.0167122701253035,-0.0126824728591692,-0.0148822347476368
"723",0.00541160652596462,0.0126165242299525,0.0094837998917876,0.017100655818346,0.00459974194053725,0.000767188235894167,0.0133737801421754,0.0189471304808817,0.0141391647180407,-0.000839266802493133
"724",0.0145042798503212,0.0174437260592211,0.00939429563434624,0.0250971695176514,0.0117118706144332,0.00536801816874877,0.0226904106532941,0.00929708276509644,0.0172225171719067,0.0289794580824827
"725",0.00116905877827533,-0.00612306352456971,-0.0113749976905351,-0.00356541617440875,0.00536746111713882,0.0021789767167304,-0.014262945222695,-0.00623157479732894,0.00304581213954513,0.00489801833895021
"726",-0.000628803072469486,0.000739306662088213,-0.0104603984464255,-0.00787230175008147,-0.00586182812322089,-0.00249992880576622,0.0165364754685042,-0.00736080422703589,0.00250066086897682,0.000812252937989699
"727",-0.0130311439255103,-0.0177298423411204,-0.0232558979626603,-0.0185140810352052,0.00178951173527064,0.00119891000111649,-0.0198822451614034,-0.0192254726709368,0.000445461024498828,-0.0142044773407461
"728",-0.00355148639828362,-0.0127848858184914,0.00757598614538879,-0.00416452541713463,-0.000210599379434684,-0.00010961261143505,-0.00760761615163486,-0.00588076727789288,0.00569901142389106,-0.00123505925958234
"729",0.0127020383024528,0.0210764143261994,0.010741096817146,0.020910296248895,-0.00126085529463793,-0.00141548643892986,0.0113823124983659,0.00957751201531498,0.0119532404470826,0.00453423541191289
"730",0.00153435263887425,0,-0.012752354782493,-0.00554207783254967,0.00631623554661198,0.005124853634634,-0.014699251686227,-0.00809140213345405,0.00384987309607254,-0.0114896742436308
"731",0.00351396966105644,0.0126834853959825,0.0172228566376398,0.0116307270028895,0.00460191307591873,0.00336289670456735,0.00396269717958808,0.00759482543675039,0.0164734589957258,0.0240763949254048
"732",-0.0162508783755472,-0.0348723488662068,-0.0084657529397143,-0.038802244698672,0.00374820140028054,0.00454152128652296,-0.0283259409425279,-0.0304300190963304,-0.0133768218133213,-0.0113497883869876
"733",0.00337667749894077,0.000763562283196517,0.0202776063893466,0.00971812072766043,0.00238638017444437,0.00161374427872918,0.0375151094122361,0.0129570326426467,0.00504085703182455,0.0110701708064096
"734",0.0123706370990178,0.021865801749646,0.0345188539369987,0.0286279986762916,-0.0111398164860764,-0.00551345705440365,0.0128971201447994,0.0264356230563372,0.0150466794798225,0.00729925362220607
"735",-0.00044947660639072,0.00273737331179791,-0.00404461902026942,0.00407835353606956,0.00083959226255681,-0.00205749352171747,0.0147795145052412,0.00138471810012808,0.0153348359686873,-0.00684387248095841
"736",-0.00782020235958714,-0.00719611344957127,0.0142132597624975,-0.00931892971635417,-0.0103848114096621,-0.00466644700149543,-0.00851469622718815,-0.0094027003021202,-0.00402754656821624,-0.000810606791958768
"737",0.00570769987871333,-0.000249946414079383,0,0.00916542179815827,-0.0105993116286393,-0.00741403243074046,0.026892784147057,-0.00111658054571173,-0.0417017449461267,-0.00811360440726594
"738",-0.0015317260762242,-0.00599990189480215,-0.00800781514315418,-0.00860419573970439,0.00128459833078742,0.0027461772292614,-0.0173856514579809,-0.00475153451067301,-0.00562636483516488,-0.00899800029003262
"739",-0.0110967111518535,-0.0223844386027588,0.00302690325234733,-0.0185629349301446,0.00149831040202009,0.00350556095087695,-0.00604685706010455,-0.0235885177020387,-0.0190964899735082,-0.00990506872576724
"740",0.00374053169604971,-0.00128645623284251,0.00301825127799105,0.00614084510886403,-0.00459368010069761,-0.00196539771585647,-0.00135204226280794,0.0115039347319714,-0.000991446624374337,-0.0125052544077175
"741",0.00563537262767522,0.00154590019657763,-0.00802399926637165,0.00585959319036156,-0.0114851217928537,-0.0033902143862945,-0.00293335678779039,-0.00625536496835288,-0.000180404192724803,-0.00548755975720583
"742",0.00424782832395665,0.00360052306056513,0.0060667769807039,0.00364061268109039,-0.000107633746170621,-0.00493905067901523,0.0144832812757933,-0.00457776152109279,-0.0135354629128316,0.00509348414873867
"743",0.00684022060342482,0.0112761036355218,0.00100513261450907,0.00677150116510372,0.00119393284898095,0,0.0194063674638214,0.00919794129661811,0.00841564215148205,0.00548978970308478
"744",-0.00464823216661914,-0.0114037309559883,-0.00803250514852838,-0.0103289652630559,-0.00444670490398558,-0.00319832209447102,-0.00919020082322608,-0.00882942382109908,-0.000272124460669931,-0.00461984469599885
"745",0.00152704896397537,0.0110227819101898,0.0151821150510436,0.00582512126334889,-0.00119851593125797,0,0.00596285713654776,0.00373593015168594,0.0125215226614783,0.01729955854448
"746",-0.0120161666398868,-0.0268762443201803,-0.0139578300320635,-0.028716132581006,0.016470696922243,0.00885283257913216,-0.00636658351219976,-0.0160323487157311,-0.0380858513517646,-0.0153464185073455
"747",0.00565734322428457,0.000260778297757724,-0.0020222488902546,0.00273274603897855,-0.00429252089834942,-0.00493611253189619,0.00773333161056033,-0.00212822157934023,0.0149990782559746,0.00421237281712639
"748",0.0101622427101236,0.00763784114682209,-0.00303938333021825,-0.00123873222470405,-0.0177819143431007,-0.0102500748426039,0.0120583238624237,0.00207335958079025,-0.0183570450213046,-0.00964764890606939
"749",0.00359327517108943,0.00833544467507896,0.00799806639215794,0.0100779809945974,-0.00559568862180526,-0.00445457704202379,0.0106156008043097,-0.00443373581209583,-0.00729311848414538,0.00720032777982405
"750",0.0019684870800476,0.0105916345952142,0.00305193152392036,0.00990337545538211,0.000220257047555128,-0.000447089029627423,0.011289205033612,0.0142519271962041,0.00357921265101657,0.0176619629297825
"751",0.00473492331355807,0.00255632008582252,0.00709947621830942,0.0100517584958086,-0.0103694679099817,-0.00358095018919435,0.0126422393223766,0.0014634419925037,0.0169873106432479,0.00578508727199134
"752",0.00213342808402417,0.00484431169512023,-0.00402814254730066,0.00339793610289552,-0.00278644353485324,-0.00269580118213497,0.00359669771679849,0.00555394758672945,0.00175343298492603,0.017666362905564
"753",-0.00141964751049484,-0.0012683534661635,0.00404443410439637,-0.00358082071136978,0.00659587203189282,0.00264058820572277,-0.0143367481283163,0.00784875557876985,-0.00994935025473931,-0.00201862644316708
"754",-0.000355206425890375,-0.00152469776290787,-0.0110777809374378,0.00437106944534205,0.00657541923507043,0.00180014837675402,0.00171174122591555,0.00490323417619609,-0.00502466730227336,-0.00121349249101033
"755",-0.00959820530643496,-0.00865128121471781,-0.00814640956367829,0.00338495857604371,-0.00476095428198364,-0.00483060430655335,-0.0194324153345657,0.00143529063504744,0.00355370803329258,-0.0028351171688914
"756",0.0169597725911224,0.0266937642497564,0.0256670934638179,0.0291568306091881,-0.000889699345979489,0.00248355470018491,-0.00239514965956455,0.0214962448953113,0.0232038490952167,0.0251827673620635
"757",0.0026472810986915,0.0010002594933376,0.00600607450208823,0.00725790752545952,0.00645784182324816,0.00439058066993203,0.00240090017480088,0.0103816731612201,-0.000910801432309705,0.00118857325538912
"758",0.000703898163194383,0.00124863707224621,0.00398028257263028,0.00209207237382292,-0.0133866656767947,-0.0040353775298978,-0.000435588572004431,-0.00527642601035316,0.0164995902415568,0.0178076370356166
"759",0.00422169842236442,-0.00324252442372541,-0.00891983671129293,-0.00579917016372289,0.00168177115268886,0,0.00893211829113993,-0.00669983668920016,-0.00618780367343197,-0.0124417099344923
"760",0.00332728722994902,0.0080078465505331,0.0120001352328758,0.0079326160890012,-0.000447184207088336,0.00123876202684992,-0.00669392518449496,0.00533953857256031,0.00496303013896404,-0.000787390854466552
"761",0.00139689780135099,0.00819263373419399,0.00889330627555163,-0.00208309499197801,-0.00548752581861511,0.000673148689152692,0.00478311012315658,0.00419342095330921,0.0132889912914882,-0.00315212641401641
"762",-0.00932644000780936,-0.0137893213378195,0.00685587174959101,-0.0160058235103083,0.0171168201695944,0.00719014357987691,-0.0168762280239765,-0.0105787483516736,-0.0209127163653118,-0.0213438275954736
"763",0.00844603749418971,0.0114855441216568,0.00583643930674449,0.00306479264107362,-0.011625753249542,-0.00479549122392897,0.0187063910231857,0.00815974177082168,0.00950314977831757,0.000807826564948932
"764",0.00270454366570605,0.000493374879024122,0.0145067484022727,-0.00258529004336971,0.0140030317294955,0.00470601737602516,-0.00345653060979345,-0.000279096524820943,0.00439302488440885,-0.0052461774260445
"765",-0.0112238933589777,-0.0180114494471931,-0.00190641065736663,-0.0115454125826281,0.00618608859073944,0.0044629518411694,-0.00910457980855528,-0.0117252265674295,-0.0104436134110829,-0.0113589960663488
"766",0.0124954955075289,0.010553066191141,-0.000955011813011386,0.0202617018839801,-0.00285490293616697,-0.00177771319830045,0.0199080005983168,0.0155367663850481,0.00595341867261934,0.00656544367339817
"767",-0.0101685819172561,-0.0256091455792955,-0.0219886830122401,-0.024065264308237,0.0101301569834309,0.00344862482894581,-0.0102962875472584,-0.0255912684617307,-0.0231348194889208,-0.0187525843160991
"768",-0.0192290219439086,-0.0308753742310105,0.00488763597752406,-0.0301650955804291,0.00457767395491371,0.00365887596123415,-0.0283916387525427,-0.019126160959933,-0.0144115932731488,-0.0124636054323451
"769",-0.0222917822117793,-0.0234331720648521,-0.0107003024915769,-0.0222167573851262,-0.00173513094194711,0.000883625870107707,-0.0229757690377653,-0.0189174471508874,-0.00186276422102727,-0.010517487817516
"770",0.00512742388592646,0.0175247438485653,0.00786625413694542,0.00732137749542194,-0.00456552887464345,-0.00220704534458405,0.00730603122689755,0.0201722166439404,0.00289264725002591,0.00467680669095438
"771",-0.0041906867662943,-0.00370955183818589,-0.0107313878443107,-0.0208020497892852,0.000327879256757369,0.00199032605294702,-0.00861288130987159,-0.0136672670453735,0.000744277984435771,-0.0110028558895792
"772",0.00475724109018638,0.0050532855590939,-0.00591757565998585,-0.0025592690070072,-0.000545680804036719,-0.00231767870302846,0.00914510855676798,-0.00353758832093853,-0.00957604145734536,-0.0145486749141351
"773",-0.0114720543132252,-0.0254038344958779,-0.00992053077216604,-0.0069283828690152,-0.000546436807191353,-0.000332089672742342,-0.00951525174619339,-0.00562131815315203,-0.000469313812722416,-0.00347368256874803
"774",-0.0108686691118034,-0.0119465966143574,-0.0140278954605488,-0.0108530857915798,0.00874216564381425,0.00387424432120875,-0.00663334328838761,-0.00684311493234557,-0.00488358363400876,-0.0113289556147773
"775",0.0155507095366327,0.0200604142154608,0.0101624922124774,0.0269073477679365,-0.00907778113151059,-0.00342983054904111,0.0181904580812566,0.0161771294970137,0.0225556721645497,0.0242397840215776
"776",0.0121033983688683,0.0161637985326653,0.0191144873935758,0.00814048670402889,0.00285270989543251,0.00166540765245315,0.0165084061448324,0.0232904823634725,0.00719888338161301,0.0215144674378465
"777",-0.00498278824298004,-0.00954407726112994,-0.00987147706269798,-0.00580394488280833,-0.011596454532288,-0.00476516642153324,-0.0115684279324063,-0.0149810556693377,-0.00394025485036897,-0.0122155473463933
"778",-0.0308658559410551,-0.0455033283478756,-0.0189430604855717,-0.045177598445246,0.0158272421580703,0.00823959553576747,-0.0373626186057852,-0.0266162969411787,-0.0398343525253271,-0.0332622435452573
"779",0.00206730183370096,-0.0190688045637842,-0.00203288489381437,-0.0111640271058711,0.00217986876455267,0.00320257630083631,0.0187050006771856,0.00120187263797766,0.00297017333610694,-0.0127923788437495
"780",-0.00721943353546606,-0.0111490431981688,-0.007128184000744,-0.00994639610936143,0.00130411777672412,-0.000879895089347271,-0.022721903432091,-0.023709551319519,-0.00611386129155522,0.000446913439102747
"781",0.0125598602287562,0.0361373259414051,0.00615391543841004,0.0325818323003275,-0.0099884787113792,-0.00539965664976483,-0.00305338083928552,0.023055763247283,0.0131680410114567,0.0178651962283896
"782",-0.00195824677413792,-0.0053012469055469,0,-0.00262922426195766,-0.0095419257585716,-0.00276946699980263,0.000707004413649237,-0.00120176503489466,-0.00275117151119741,0.00394900110499585
"783",0.0104663157373366,0.00729310949508344,0.00509680109341626,0.0263640619807803,-0.00542615094844923,-0.00122222069168243,0.00870946796316874,0.00721996633250011,0.0191209469428955,0.0118007183910438
"784",-0.000832662077561275,-0.00863273928529207,-0.00608526102565454,-0.0125865948967366,0.0041194640367932,0.00233605834855344,0.00910183416506904,-0.0062720986670286,-0.000840063497808186,-0.00561547411050289
"785",0.0157354054164858,0.0230339076249522,0.0102039746030314,0.0257544715836457,0.00188505784101745,0.00221962371503914,0.0268269157381149,0.0135253570441207,0.0241031574728778,0.0304082808699191
"786",0.00473824673929868,-0.00109843127581333,0,0.00355086690838524,-0.0113983560582998,-0.00531531552684994,0.00945994029262698,0.00207592539837242,-0.00337532375364014,-0.00505895277612167
"787",0.00589517325087385,0.00494786589263407,0.00202023505990989,0.0037904737138077,-0.0040303757509057,-0.00356181286927137,0.0133864610096497,0.00562308774108899,0.00668194965675051,0.0088981828450192
"788",0.00207368241103989,-0.000546980888919468,-0.0161290259786369,-0.0085597800044992,0.00539549973463016,0.000559242029515294,-0.000219894884041949,-0.00971151679145565,-0.00463722482349815,0.00588001847142516
"789",0.000180124226383693,0.00136846404306357,0.0122952521261634,0.00126954508651367,-0.00413662098895207,-0.000781966413007096,0.00418380641429628,0.00267459863993214,-0.00365397822550495,-0.00542802922543661
"790",-0.0121449133360039,-0.0210444262158427,-0.00404840781499427,-0.0230787930367874,0.0156039453658734,0.00759786090508352,-0.00789469645007179,-0.00859516256301351,-0.0108187494269734,-0.0163728741687471
"791",0.00919772237076533,0.00949246679558091,0.00203231125513792,0.00960536103255638,0.00243120523832641,0.000554927579841324,0.00972616164118878,0.00956638272146959,-0.00491239229689866,0.00810937083926322
"792",-0.00135328335663221,-0.00885002364131282,0.00202843038530998,-0.00822837045127622,0.00562389135594077,0.00365685454846365,0.00503437200243217,-0.00444193101865697,0.00884870520819003,-0.0169348735900949
"793",0.000632223895218997,0.00502260750839922,0.00607294248459023,0.010111431506026,0.00515349877743021,0.00154598240391901,-0.00239573773032786,0.00832861383520056,0.010340707420196,0.0176571726432413
"794",0.0103849148510506,0.00222076213499212,0.0100600457354689,0.0169406339568599,-0.000437940900656297,0.00103897156353305,0.0102625972093067,0.00855485985442006,0,-0.010156572821003
"795",0.00277059769140142,0.0132963428390889,0.00298830392225602,0.0113579253688145,-0.0013132506930188,0.00055316566432273,0.000432034352852995,0.0152089010628293,0.0145298090103263,0.0106884025606933
"796",0.000891036819194335,0.012028581291982,0.00695165930691699,0.00124787115362368,-0.0025223920841343,-0.000993829419531522,-0.00216085776145691,-0.00316938195452754,0.00549450564297893,0.00972926960187404
"797",0.00302793386987998,0.00135083215383935,-0.00986249914082837,-0.0052344456837311,0.00527547125568484,0.00176699389508972,0.00411396903541417,-0.00115591752719657,-0.00716648769595518,-0.00879774891871954
"798",0.0142933063193504,0.0207712649064384,0.00996073689994614,0.0260586060660462,-0.0131183721857153,-0.00474162644793452,0.0228545386837922,0.0205438835302951,-0.000180492643138241,0.0118343758967849
"799",0.00017481809057629,-0.00396424212392943,0.0069031106964037,0.000732761438573037,-0.00520646709803285,-0.00266027529627033,0.0124369467125063,-0.00481992348757276,-0.00839275351308999,-0.00125311570013642
"800",0.00166255577157415,-0.00159170876804759,-0.00391779064354991,0.005612074194145,0.000222314264102241,0.00255653201345907,0.00333096638247432,-0.00113924731221204,-0.00145609760073084,-0.0108741776279682
"801",0.00445602697554293,0.00425200574462226,-0.00688295411242212,0.00703760894427807,-0.00256114045224931,-0.00166339535647742,0.00539560061122879,-0.00912753975660319,-0.011392635696385,0.00295987758725458
"802",0.00417511659985226,0.00846753241649245,0.00990088467347916,0.000240533903196116,0.00368390465391966,-0.00088809472019602,0.00495355428052591,0.00690843091015014,0.00119846039274951,-0.00252956316850506
"803",0.0000863226856009369,0.0047235113251618,0.00980381820011988,-0.00337260736952938,0.00622755461858926,0.0015562695271536,0.00739355238866968,0.000571808114484984,-0.00598527635332002,-0.00591707919774553
"804",0.000259797002732043,-0.010707918729845,-0.00485421729542601,-0.00725167970656837,-0.00132608958875902,0,-0.00285430373508511,0.00171459748320046,0.00379809181467605,-0.0119047301272583
"805",0.00796634593102863,0.0163674549265582,0.0097560231926479,0.0129047944763818,0.00796783139535795,0.0038829651097656,0.0259659501819682,0.0168280811140986,0.0188261441599655,0.0133390202979642
"806",0.00592719660934149,0.00285730338639834,0.00386456734590435,0.0108176960234461,0.00428185785924651,0.00121584562302313,0.0121563089693435,-0.00112207290324784,-0.00733701073664839,0.00891716287918798
"807",-0.00051224258829774,-0.0069931721252432,-0.00673690024300311,-0.00761004794804854,-0.00327963712362356,-0.00264897588413271,-0.00393792682390648,-0.00224671701160439,0.00684369036750399,-0.00210443502469138
"808",-0.00506177865351509,-0.0112151840973744,-0.001938245868777,-0.0129407070348394,0.000986863227195656,-0.00132841885868207,-0.00849949666626559,-0.016198899314217,-0.0186695402816581,-0.01223100333295
"809",0.00534610723154771,0.00131871987319632,0.00485444804070578,0.00364185233729719,0.00109666083783644,0.00332421703109187,0.0103667558661935,0.00660946455038824,-0.00489470820922344,0
"810",0.00703315274488747,0.00579571843180093,0.00966184892204258,0.00701514347292953,-0.00470722488116671,-0.00209907292777867,-0.00276217695729375,-0.002569381205621,0.00529002320185601,-0.00426988417232754
"811",-0.00485484291746063,-0.0154532222556109,-0.0162679503371341,-0.0148932434125751,-0.0182550094215829,-0.00996093063370151,0.00316586476700143,-0.0151683545109769,-0.0186484213441653,-0.0111492962624892
"812",-0.00162604147071743,0.000531993119428753,-0.00583641040747196,-0.0026821588757705,-0.00638499144176063,-0.00368857057469063,0.00157332533215482,-0.000872496197010575,0.00451548435045668,-0.0056373907344931
"813",-0.000600115166536241,0.00771078589349528,0.0156555378202778,0.00489000698847986,0.0028177308837769,0.00235585444221953,-0.00357943829821616,0.0116348343811705,0.0169507119025165,0.0017444157174622
"814",0.00634757129355434,0.00949860321168416,0.0125237996727834,0.0180046706195074,-0.00382233397644249,-0.00145466925208937,0.00439048283225962,0.0212767931259361,0.00147346906615597,0.0226382280421098
"815",0.000681856722046792,-0.00444325786002253,0.00570905521679932,0.00382400325559673,0.00315997803814416,0.00100815849482849,-0.00198696374834428,-0.00281557961077317,-0.00717240459770119,0.0021286238789695
"816",-0.00340704498648647,0.00656334422344118,-0.0122990175524946,0.0028573229286204,0.00686225699688281,0.00235169127270862,-0.00895894627678806,-0.0095989332963996,0.00907655821916675,-0.000849649729898538
"817",0.00683737466163392,0.0164321602110333,0.0153256345187631,0.0261160588936162,-0.00244509633666057,-0.00207180920739036,0.00462034606513373,0.0193841349213275,0.0120239103815671,0.0195577740490089
"818",0.00814965686078839,0.00538850715993378,-0.00283009455135741,0.00902334707581476,-0.0166376344736844,-0.00898324549285245,0.0207960301215795,0.00531316571907681,0.00571374014667625,0.0158465370998924
"819",0.00235763435185943,-0.00689111918667551,0.00283812671831907,0.00298104750467321,0.0016001916960402,0.00294588958303188,0.0201764281726833,-0.000556251682812592,0.00126251241106057,-0.000821006858102935
"820",-0.00571259083277875,-0.0110513840568808,0,-0.00868760171591243,0.0127842143656007,0.00621329715328778,-0.0215058108946936,-0.0158641792045926,0.0131495903192793,-0.00369756658899045
"821",0.00346431344575571,-0.000519545867308957,0.000943103266584755,0.00345915731075586,0.00045026767227796,-0.00112279060459408,0.000392217925669902,0.00735308833793646,0.00142238423721897,-0.00164954680753537
"822",0.00656721042535247,0.0145606028577647,0.00282798800349338,0.00620562337097486,0.0023662840890244,0.00112405268038263,0.0158893415965913,0.0106678446594868,0.00878825550309359,0.00206531912904606
"823",0.00158925422647971,0.0079446855992058,-0.00187972947888937,-0.00799429810179353,0.00528141907378621,0.00269424060177537,-0.00656525669002683,-0.000555231578312054,-0.0055437962473055,-0.000824475860280893
"824",0.000751689106683884,0.000508317306082029,-0.00188338141234645,-0.00207263900849164,0.00324236131822664,0.00190316516503186,0.0227405603759572,0.000555540031680568,-0.00283160777220404,0.00371290560147886
"825",0.0113492284677508,0.0142311400987685,0.00471716991665949,0.0147670794012642,-0.00702029852445807,-0.00268156433256006,0.000950119126654325,0.0127779518842543,0.00301709995532695,0.011508480076293
"826",0.000825062692280554,-0.00350778659158801,0.00469466005850383,-0.0054570270861235,0.00112204870021304,0.00168044927940314,-0.0248717860634572,0.000548421936290566,0.00548529598766079,0.00365708345691451
"827",-0.0159120047865183,-0.02137287976066,-0.0186913926142843,-0.0292636089986644,0.00728634296451336,0.00604059254206257,-0.0208331484957525,-0.0216555570741785,-0.0212054901679632,-0.0182186646443475
"828",0.00376998521473659,-0.00385434378106442,-0.00190499051833692,-0.00400393776184693,-0.00244842271539436,-0.00244576876912528,0.00377792376995001,-0.0050434842371202,-0.000809025544930342,-0.0127835421184697
"829",0.00893058739887387,0.00851193317151533,-0.00381674260748488,0.0118232907202811,0.0035699664262796,0.000446080988985686,0.0156498868333403,0.00816654326659028,0.0027889968009176,0.00793648541716063
"830",-0.00181952460349266,-0.00818401585341799,0.00383136594513256,-0.00327171929412207,0.00822587692060606,0.00323117647600357,0.0187243747224559,0.00139675479451995,0.00762604528643496,0.0049731226595251
"831",0.00298349126344988,-0.0108301726978757,-0.00858789764893308,0.00422020742037921,-0.00297693666810062,-0.00233229093749432,0.0145508509220105,-0.00223141209262667,-0.00418486339924962,0.00247419288560891
"832",0.00652760652427498,0.00860233286580425,0.0067375292959988,0.00537010484253742,-0.00353833473331233,-0.00278313156804499,0.013021342851226,0.00698918118647152,0.0120708695304317,0.00658156363703033
"833",-0.00377650389267659,-0.00155035558053362,0.00669204116614019,0,0.00110926960924584,0.000669988597674198,0.00633380071260747,-0.00111044014664263,-0.0038872867941111,-0.00490381329421719
"834",-0.0236502240521478,-0.0445251980360979,-0.0180438081462552,-0.0357641254606517,0.0140783213377988,0.0093712351089521,-0.0316545711756765,-0.0330740284713151,0.0166740310421287,-0.0151951590075315
"835",0.00759612949867994,-0.00487678112699297,-0.00386842027007395,0.00842953046851225,-0.00852625453582334,-0.00508471501693042,0.00344101581896861,0.0063235538482278,-0.00279158168345772,0.00333606789495611
"836",0.0123973844415497,0.0185136367865357,0.0116509637292936,0.0164795171685599,0.00418970694991749,0.00166631618409885,0.041341039148258,0.0159956724636672,-0.000262435487051516,0.00789703081839277
"837",-0.0169617487315843,-0.0155040908253133,-0.00287963744982189,-0.0119827706629595,0.0115278754344568,0.00609982255767072,-0.0311014210303145,-0.00590403991908561,0.00945049010719701,0.00783502902155764
"838",0.0129617989739328,0.00705981927149435,0.00288795370947703,0.00546950793545875,-0.0013068101828706,-0.00262051363806759,0.0309664865977444,0.0152717600764867,0.00320736821075451,0.00490995854541798
"839",-0.023514549992082,-0.0401728130034278,-0.0307104306021803,-0.04588445523878,0.017995441105249,0.00676205417974107,-0.0234428912911945,-0.0406686241204169,-0.0074310894124836,-0.0268729322961048
"840",-0.00595676672247414,-0.0269662565448211,-0.00099011494022283,-0.0180963623332494,0.00589200487881758,0.00385346501682382,-0.0140658807161048,-0.015389186958487,0.0019151475080923,-0.0225941773588147
"841",-0.0332132657261301,-0.0534063138491681,-0.00594645966266871,-0.0408985681268305,0.030887331143473,0.0109680785263109,-0.0401372004542252,-0.055145896708145,0.0295421158933744,-0.0196918202787819
"842",-0.0148752922575006,-0.00579455693791331,-0.0089730769777594,0.00526404920381385,-0.0125008956988562,-0.00271168077508621,-0.0168451670384201,0.00530574845609255,-0.00185670523852988,-0.00524014825566066
"843",0.0440411026205816,0.0763805688940289,0.0281690486027826,0.0720086564121503,-0.020716362762176,-0.00761553638100476,0.0659141187510042,0.0509158824216644,-0.0059186354760794,0.0193151962987981
"844",-0.00284092815223191,-0.0054147479930714,-0.0225051953446688,-0.0180750690809538,-0.00256341060652188,0.00120611147826222,0.00113466077378854,-0.014180149854548,0.0262822488730119,-0.00172262936785217
"845",0.0139858143998659,0.0163322873031591,0.00900912662222964,0.0124376411805602,-0.0076049228026448,-0.00251862093413524,0.0162451599774593,0.0107881425304912,0.00613291874248567,0.00819678682120339
"846",-0.0124303779829975,-0.021990359280469,-0.00793648945761061,-0.00933662744814268,0.0065841285075523,0.00274437095688329,-0.0131972475239297,-0.0103765166926297,-0.00691930795849582,-0.00855803888595574
"847",-0.0181052205080607,-0.0302683343944699,-0.00699987587808526,-0.0205852073955258,0.0173705938138713,0.00645845829186031,-0.0308909691720481,-0.0170756098313831,-0.00157593731877792,-0.0254639689982534
"848",0.000526674349315082,-0.000594296252144244,-0.00201401143790236,-0.00607748917604789,-0.00368886564154114,-0.00217509900829194,-0.00155479520778967,-0.000305286293781126,-0.00839081145491039,-0.0283436440301731
"849",-0.0136023996896749,-0.0190365604004807,-0.0171544842501318,-0.0208916760578096,0.0153387245205541,0.00730337261949954,-0.0255013176846196,-0.0216464026873832,0.00108911694797986,-0.00136734681240436
"850",-0.00569395606258161,0.00424524393786618,0.00718682155159489,-0.00962814887964136,0.00333445663062037,0.000865228773265558,-0.00839022905710196,-0.00218156446925188,-0.0239350660964945,-0.00912836160459607
"851",-0.037759537023286,-0.0314009287748945,-0.0152903729964058,-0.0496582817511254,0.0210789991731086,0.00973097214158325,-0.0483477006897396,-0.0371640053426897,-0.006773566152111,-0.0207277302351985
"852",0.0145992741122376,0.0199502815097747,0.00931655013226407,0.0323471793284136,0.00101725654755014,0.000535338534906282,0.03238735131791,0.0204347748155094,-0.00535216696658036,0.010348075457902
"853",-0.0128312985461553,-0.0259782642729364,-0.0133335189984637,-0.0104443739787277,-0.00345375040865059,0,-0.0200941654169773,-0.0171647227264558,0.0140600155002604,-0.000931085981564328
"854",0.00102153636888724,-0.00156881663037101,-0.00623695410361369,-0.0108254072714297,0.00489309343475886,0.00342477820838871,0.010462289734398,-0.00840884846886669,0.00445057358612022,-0.00792165449983961
"855",-0.00602876200204261,-0.0141422266199784,-0.0125525996608388,-0.000547521130797368,-0.00284003388147636,-0.00202699987686772,-0.00393393260384478,-0.00913220823504579,0.00945807762902118,0.0108030940099144
"856",0.0334983321754494,0.0621613764154167,0.024364875341675,0.0604984431385753,-0.0226882871567041,-0.00951064933905832,0.054261472306901,0.0513495266596544,0.00185701863883669,0.0292750765132741
"857",-0.0125495897567045,-0.0204082163285458,-0.0165458871152572,-0.0165202018984233,0.00458056061484857,0.00453141893763864,-0.0149868893256772,-0.0159677474985794,0.00160076667620235,-0.00857780778638462
"858",-0.0168238547948674,-0.0119482488595812,-0.00315449982860627,-0.018372851605969,0.00702812915012951,0.00129263522085976,-0.0194195035924216,-0.0104993819589173,0.00866425829401729,-0.0186703822178462
"859",0.0260393997823063,0.0310076448403775,0.0052740951945085,0.0350267187213851,-0.00949828441030798,-0.00570106758355038,0.022049733457018,0.0369773260881303,-0.00108418810493904,0.012065039772875
"860",0.00344397143220676,-0.00210526106821263,-0.00209854508085894,-0.00361671806820607,-0.00729686255896844,-0.00140669715738184,-0.00259702931323202,-0.00279081105147905,-0.015194523419557,0.00550208235748162
"861",-0.0351367956624009,-0.0491259839275837,-0.0189275612766411,-0.0355195432854208,0.0268816725328909,0.0138677136594534,-0.0542756845227046,-0.0407334394802956,0.0104272889998924,-0.0310077024594181
"862",-0.0124505964547102,-0.00919184341254553,-0.016077143900191,-0.0155914814746622,0.00766954698773281,0.00406070777231005,-0.00508253764265831,-0.00842810117465742,0.0192968869989614,0.00188232704909397
"863",0.0107118561359958,0.0111965389876387,0.00980375626786012,0.0229380811078681,-0.00497249539104572,-0.00308645022059861,0.0174543110842913,0.0117686212135992,-0.00403323736987793,0.00798490818368358
"864",-0.00534598148512555,-0.00284712275503851,0.00107879829651014,-0.0053388625033991,-0.00112183489321249,0.000106697072237649,0.0050204623611112,0.00387720552529869,-0.00363638016528933,0.0046598644724829
"865",0.0292313543647078,0.0491751225158119,0.0172409874219273,0.0348898813429483,-0.0178677681372251,-0.00928671077869092,0.0418402082328861,0.0379786321677353,-0.0131884292167954,0.0166975025710112
"866",0.00485595983056841,0.00332617294918358,-0.00211811286415886,0.00518649552402617,0.0126829926064596,0.00635725922194497,0.0103898674348466,0.00186054070098596,0.00874170792013351,0.00136868840960847
"867",-0.00154997642821142,0.00693185017966225,0.0063695609371861,0.000258119180829741,-0.00513308066023688,-0.00085638713864733,0.0118639984007147,0.00185736137720061,-0.00341641524178959,0.00273344776777806
"868",0.022737297918793,0.0359174437786274,0.0179321179570693,0.0301777788442947,-0.00412744627384898,-0.00310831653631372,0.0216929790216087,0.0299653502095947,0.0116220737729444,0.0168104514110876
"869",-0.000356868073041361,-0.00953479554113368,0.00414548412684868,0,0.00569920258865175,0.00279502550557731,-0.00726858134307562,-0.00419895742795162,-0.00545496331027306,0.00223419928982249
"870",0.00160749228105317,0.00554245290587851,-0.00206423100550435,-0.00500738813987545,0.00813884382151175,0.00471638549039555,0.00154142866225082,0.000301485526305267,0.0130474526211677,0.000445917171275401
"871",0.00108436114701216,0.00116037132839986,0.00206850086913324,0.00452958465620967,-0.00163537931374136,-0.00202660482206074,-0.0028855378477558,-0.00671323728568096,0.00762920414062007,-0.00178259847966811
"872",-0.00286413044252087,-0.00663019222799577,0.00722356683506264,0.0172845959161263,-0.00286580546988746,-0.000748576503408316,-0.00713895649513852,0.00214055776306821,-0.0198648779636101,-0.00401780231396276
"873",-0.0165154536740671,-0.00923706197976371,-0.0122948868582701,-0.0192073262104436,0.0119083949290952,0.00599111895374094,-0.0281772998956471,-0.00762879719008247,0.00880470146029322,-0.00224111676075323
"874",-0.00310316081721929,0.00661634116503618,-0.00428393375989622,0.0025779631635745,0.00679719195565487,0.00372253974196246,0.000599947983138671,0.00492008749816897,-0.0041169206451277,-0.0166218384377776
"875",-0.0165703787261433,-0.0179265036998895,-0.00314775702001047,-0.0176454500460691,-0.0059451056430051,-0.000848095925587433,-0.0205999531043317,-0.0140758950371839,0.00289380743018963,0.00228421090344666
"876",0.00418907621324172,0.0021296454319335,0.00421051062826971,0.0118038568665089,0.00405442951759372,0.00159074485234711,0.0255196715213581,0.0117938780119384,0.0120362651598616,0.0182315253844831
"877",-0.0031521459072491,-0.00394637642736384,-0.011530386461215,-0.00684737338794916,0.00938943922458391,0.00709423807892695,-0.011438702345225,-0.00797532577350879,-0.0136038283870344,-0.0107431451285394
"878",-0.0308750775593342,-0.0374887143732396,-0.0243903095113993,-0.0406028213123525,0.0109022239582441,0.00430956474747202,-0.0320748001535045,-0.0281385420944603,0.00148650595380317,-0.0276017606022768
"879",-0.00949973063485687,-0.00728325857006673,0,-0.00665430388078225,0.00672802720240284,0.00146585032766056,-0.00985726292668165,-0.00827226712789064,0.00338091044893818,0.00372261089084946
"880",-0.00445679304306734,0.0169062024779028,0.00326076146503618,0.00723461069916298,0.00157678673418049,-0.000440453518088413,-0.00190646183363841,0.0134742780326778,-0.0381327991452992,-0.0152989615223466
"881",-0.00544974742403437,-0.00470514390695842,0.00433367910220239,0.00425661507520303,-0.00797228182484766,-0.00178249204044478,-0.0191000655751877,-0.00158271828705281,0.0123889011244966,-0.00188311652441298
"882",0.00655609481093866,0.0226915167244539,0.0204965338126992,0.0185429788399543,0.00823534580228946,0.00241618304608737,-0.0194717906693911,0.0117310962882409,-0.0167102374328676,0.00283005256186408
"883",0.0314960140956468,0.0354389524589309,0.0190272552744088,0.0221064720830657,-0.0117107159027462,-0.00314370408642861,0.0476606477842461,0.0363522880365899,0.0104712125916879,0.0225775443640059
"884",0.00989542553742062,0.0104167205059817,0.00207480369529844,0.0048348137992138,-0.00637220237252056,-0.00241706832177679,0.0107413237253755,0.000302387870286802,-0.00441691995879756,0.00919974372801868
"885",0.00746568333811215,0.00147272759500128,-0.00621094324897198,0.012155032672714,-0.00571269150445586,-0.00263407366516999,0.0131276239670333,0.00030240329691722,0.00981146668212163,0.00182312908320581
"886",0.000647965426826547,-0.00264701134435119,-0.00520865066279996,-0.00800587544018261,-0.000402352185643662,0.00169045591468908,0.00370222711125434,0.000906401604853446,-0.00861781844695997,-0.0113739613018505
"887",0.0150886114398023,0.0253612706694535,0.0052359227553298,0.0116012933333998,-0.00857023751408514,-0.00495747194528839,0.0219263691013787,0.0132850349800788,0.00869273082300093,0.0161067811886209
"888",-0.0000912037954093892,0.00258835298845361,0.00729157631658262,-0.00199460715486999,0.0100679347972632,0.00498217091784015,-0.00581516574168106,0.00327754306955175,-0.000506911114338315,-0.00181156937638549
"889",0.000273715070989944,0.0100400193523931,-0.00827322127816699,-0.00474624020723036,0.00996778205253324,0.00516740710294683,-0.00221896448264791,0.002079363129176,-0.0005917159613259,0.00952804655642714
"890",-0.0275344730453413,-0.0312409898230332,-0.025026131008871,-0.0298697450999976,0.00488488446418867,0.00577061107515364,-0.0307251491084874,-0.0222290471050116,-0.013194662610302,-0.0125843292251807
"891",0.00590624680414953,0.00586351491524661,0.00320854461086495,0.0131957449509237,-0.00615083350334444,-0.00260746903369036,0.0114701942731892,0.0142467499772352,-0.00805686994183386,-0.000910226211123244
"892",0.0110916639692507,0.00204002773609013,0.00639634543780976,0.0234932643686543,0.0014975801337771,0.00104567310677073,0.0171133748415422,0.0140468423836104,0.00794952887022737,0.00820039019244789
"893",-0.0129982178688194,-0.017161029559181,-0.0180082893867024,-0.0102296858681462,0.0169437022782621,0.00637283244628328,-0.0192581116048138,-0.0132625024920511,-0.00685815676196899,-0.00271126125667331
"894",0.0223220469377188,0.036105146112918,0.0183385350324958,0.0302494190878344,-0.0115649227367113,-0.00550195565046563,0.0359652572777365,0.028076365755644,0.00871819609353808,0.0199366670670988
"895",0.0086790433552435,0.0131392926756206,0.0148307713477767,0.0068508212296019,-0.0106098729445389,-0.00323637213829553,0.0117714773079676,0.0136545488671933,-0.00658912368142117,-0.00310973207646137
"896",0.0104157158669897,0.00733019632270726,0.0010438991537689,0.00680456957096687,-0.00170387610622336,-0.000313879220935287,0.0258336663594536,0.00917175538960269,-0.00490997518855973,-0.000891345105075714
"897",-0.0000897389234056911,0.0064372401022097,-0.00521371449830554,-0.00168926977866235,-0.0096376973039245,-0.003457351395594,-0.000192308410412401,0.00198816565909188,-0.0173995416568441,-0.0107046737841719
"898",-0.00645444163516828,-0.00834286384728167,0.0115303555431803,-0.00556101857199709,0.0032437840127777,0.00431003370471394,-0.00153881978922366,-0.00935341051800742,0.00237861858199961,0.00405774690872085
"899",-0.0048723569571264,0.00224333225614526,0.00621759377488695,0.00170183276601055,-0.000302502801797666,0.00209340757289422,-0.00885767072153454,0.00457774985039117,0.0044823519465842,0.0143690478374703
"900",-0.000181287386889495,-0.0016787991536733,-0.00823902041355917,0.00485435134438905,0.0155647087934494,0.00585010584667867,0.00349722687561016,0.00113952436823617,0.0104995799238814,0.0132802587701601
"901",0.0225807523798716,0.0369958029056761,0.0218072355396639,0.0258455367788359,-0.0140382042456888,-0.00309275118291452,0.0303971191545509,0.0301560111961632,0.000432963900475647,0.0192223290506586
"902",-0.00478879841183721,0.00135103593551111,-0.00406547431897597,-0.00470927680814792,0.00577201141047334,0.00470059759180597,-0.00526103909178932,-0.00856099738698901,0.00389472906443888,0.00342901439923127
"903",0.00668344022315215,0.0008098112776731,-0.00204071890804347,0.00141939413914649,-0.00765170673717375,-0.00415864125778787,0.00321115060930155,0.00334275486395419,0.00629367197678543,0.00854337299574337
"904",-0.00106230203349411,-0.000269282997078624,-0.00102267217371699,-0.00448835284235938,0.00466652055173311,0.00480174287161406,-0.0124271532819856,-0.000278015044209878,0.00222757023451359,-0.00465902280095076
"905",-0.00407655200320756,0.000539437379233565,0.00921205298595451,-0.00142389078385463,0.0109076521968761,0.00654567273288453,-0.00324126262784685,-0.000555301415900877,0.0073516240207312,-0.00893604810459558
"906",0.00533874743017049,0.000808610925989495,0.0010142549714649,0.00522814102681379,-0.00369703077545913,-0.000206096593837413,0.00994656273118544,0.00611278960481076,-0.00373382565287939,0.00343490326253937
"907",-0.00539858501843404,-0.00673479337512484,-0.00607900519218851,-0.0137117150392053,0.00210633385904457,0.00505824230187457,-0.00776549174800489,-0.0107703736179992,0.00281091136608325,-0.0106975486074448
"908",-0.0274069225019203,-0.0461080296802242,-0.0336389902692403,-0.0318789217861368,0.0134073727618715,0.00565023277452625,-0.0240504147046017,-0.0337799488471114,-0.00331272394514415,-0.0224913537169457
"909",-0.00613012626833442,-0.00255902986073275,-0.00316460707873734,0.00173276598795624,-0.00246828739712501,-0.00255399673631052,-0.0115390658370678,-0.00115562932757884,0.0121868165054311,-0.00752215774694576
"910",-0.00294578590978345,-0.00427578748701452,-0.00105863403654638,0.00543747440918141,0.0124718905412802,0.004301138634631,-0.00217649524894592,0.000867494740516062,-0.00025258062438116,-0.000891650799776267
"911",-0.000461611896092284,0.00601187706752571,0.00741569812956833,0.00934123368755468,0.0250263358554572,0.00723994284904927,0.000991508447125033,0.00289031747476343,0.00833758646349314,-0.00312356292659821
"912",0.0122851258059271,0.0108140769419465,0.00525754162870506,0.0104726447114809,-0.00572207383579737,-0.00506180526471522,0.0217909088060146,0.019308140661447,0.000167017451757623,0.0143241167204717
"913",0.00182525277231904,-0.000844693027592935,0.0062762816575459,-0.000723144035991052,0.00268587068452453,-0.00101812573677429,0.000193749196158999,0.00452359356503029,0.00392485177453028,-0.0039717927589521
"914",-0.0173971642112378,-0.0166244437257452,-0.002078871467322,-0.00771815832899558,0.0155939830359153,0.00448215181878808,-0.0226788979708881,-0.0115393095234081,0.00141405754937574,-0.0101905157808873
"915",-0.00324422048600315,-0.016045866051334,-0.00937517791573417,-0.00291688233867515,-0.00113059568966811,-0.00324450343810534,-0.00297505714679913,-0.00740341606021866,-0.00348864526529324,-0.00626679242697858
"916",-0.00381283074464278,0,-0.0063091554073702,-0.00902032910514206,0.000188533741477093,0.00132246630091859,-0.00477426010751014,0.0014344056102864,-0.00158374592328292,-0.00675680343109109
"917",-0.0148432326208736,-0.017181174891581,-0.00105863403654638,-0.0127916187537132,0.0160281408916481,0.00792408131729117,-0.00439736511063848,-0.00887999938447925,0.00484222745735696,-0.0113379006567939
"918",0.00388526666931721,-0.000888912892838878,-0.00317723682881355,-0.00647920916116873,-0.00324749578593431,-0.00453543383589827,0.0130499937676674,0.00780339242669714,0.00830840803997668,0.00504599179799725
"919",-0.00670181508728773,0.000296674384352658,-0.0010631024128156,-0.00627043358591239,0.00940327513789652,0.00455609771563736,-0.00554917991981829,-0.00286727903530504,-0.00329599535847069,0.0114102993379197
"920",0.0154899042317291,0.019567158678391,0.0127660047148734,0.0219588503103352,-0.0283162973722335,-0.0114908284979919,0.0159426141084666,0.0192693140121976,0.000413384593364707,0.0171480117157852
"921",-0.0145049708452017,-0.0171561940957476,-0.00315131075392272,-0.0165471178548051,0.0191743122384636,0.00764762236763183,-0.00921930486911215,-0.00846533119361137,-0.000826361444072998,-0.0017746899064317
"922",0,0.00562128068207035,-0.0115912303900673,0.00602677273080277,0.0110831457215921,0.00445253778040455,0.00930509134303859,0.0082527280286806,0.00967660211143473,-0.0133332888102071
"923",0.0299116033224947,0.0385408494474702,0.0277185765234491,0.0351972258505686,-0.0206767410141256,-0.00720085957299077,0.0315808719760116,0.0273782412879864,-0.00319462642210622,0.0198197805590823
"924",0.00931234104293277,0.00821522584377155,-0.0031118689725208,0.00168799990593382,-0.0105657894558577,-0.00417114754761327,0.0125503437773791,0.00576906524452769,0.0049305529635868,0.00706713234755285
"925",0.0129715121417449,0.00983400894649367,0.00728365257859931,0.0117954886466942,-0.0123945773271954,-0.00571983343748594,0.0131450620319595,0.0106530817393677,-0.00351623187900707,0.00526322156738601
"926",-0.0112723846699225,-0.0178071788260012,0,-0.0145130058044683,0.0204666567316043,0.00791081031362206,-0.0139014101568598,-0.0132434829944293,0.00689312319962965,0.00523562019718837
"927",0.00702290436955399,0.00736530651097844,0.00206623066081546,0.0108640498190888,-0.0079465293011004,-0.00275223610684194,0.00056379687180419,0.00520408495646185,0.0000815158944136307,0.00217010912772109
"928",0.00461913841074324,0.00899879005574222,0.00309298564034388,0.00573205475297689,-0.0197411695346346,-0.00787084462010634,-0.00751441043688861,0.00844679027217965,-0.00937169757453915,-0.00563024417114466
"929",0.00504873890151281,0.00641033000804669,0.00719406664415323,0.00356230798470492,-0.0045722163065286,-0.00288533004377323,0.00397471958898166,0.001621130454043,0.00139852749915326,0.0104531334813114
"930",0.011122845450505,0.0160620813781851,0.0102044071799308,0.0238995158736994,0.00488645418747358,0.00475323048034637,0.0156488784391506,0.014836890873192,-0.000903639179241633,0.00732757416011309
"931",-0.000620756226571539,0.00953947006327915,0.00303014250524458,-0.000462235311782466,0.00962889711159232,0.00503929339331322,-0.00297052917411722,0.000531583390435575,0.0197335466271942,0.00299525195401307
"932",0.00381718837385536,0.000539838052945552,-0.00201397251727442,0.00138734721622003,-0.0148350068167044,-0.0034794412625877,0.00781974443000344,0.00106297749658513,-0.000645016948355503,-0.00170654908078371
"933",-0.000265674312781572,-0.00215855039802149,-0.0131182510863742,-0.0050795475639227,-0.00987549235493301,-0.00349044642339869,-0.00535732655865939,-0.00371557966452207,0.00556716950835612,-0.00512813520556832
"934",0.000373434820160945,-0.0102759312071197,-0.00306741333487415,-0.00162453817937525,0.00404876373179563,0.0022661857679096,0.00297199393039094,-0.00583069285720239,-0.000722105449460941,0.00343637901994409
"935",0.01529034740573,0.0193988178011477,0.0174358336117033,0.015806634326595,0.00580266506848037,0.00308474282644666,0.0224072274149143,0.0172969416989281,0.00264976712180998,0.00813358273024756
"936",-0.00201340289512786,0.00268041539907782,-0.0110886400490582,-0.00297534932181398,0.0138867941544993,0.00932661121179845,-0.015757981583796,0.00239139080692219,0.00912948644679701,-0.0106157845556669
"937",-0.00491315146410565,0.000267411364072601,-0.0030581829590911,0.000688850382142281,0.0089699377240009,0.00152279847228476,-0.0103055347233412,0,0.00150777713661165,0.00600867863313748
"938",-0.00811150978804964,-0.0117584934104733,-0.00408996487133584,-0.00642197243859033,0.00286788430914875,0.001419843900065,-0.0224320729909921,-0.0108666172782984,0.000792440589360677,0.000853142814789987
"939",0.0206219741285871,0.0316387735254979,0.013347065338152,0.0184673544460572,-0.0134401977146948,-0.00496084645457961,0.0272447099704356,0.0262590473635027,0.00308787799474564,0.0153453669436308
"940",-0.00479015146593564,-0.00655313822116055,0.00506580777585386,-0.00181340458951296,0.0173909572144915,0.00773238808614751,-0.00989882935730146,-0.00626599139892181,0.000236790587468727,-0.00671712532960733
"941",0.00350077409962601,0.00897109917916716,0.00403224355735854,0.00726620285138058,0.00683778799571533,0.00333206051085155,0.00264079063380862,0.010509522256573,0.00891727423518573,0
"942",-0.00174423792810952,-0.00470727422802308,0.00502015117549837,0.00338151039245904,-0.00414998925550625,-0.0024154099970205,-0.00733787509678385,0.000519917665885883,0.000782158792055565,0.0131023214391592
"943",-0.00297053020192628,-0.00551775243421138,-0.0119879092532178,0.0058412054339132,-0.000663790875962023,-0.00121034519062135,0.00227453386185772,0.000260142436406596,-0.000312567416472787,0.00584064025226727
"944",0.00420585047859756,0.010568235007903,0.00202226691626861,0.0147420284636404,-0.00483198562073606,0.000536359344962989,0.00491662801935311,0.0161078411863416,0.00781799678467676,0.00207379995796053
"945",-0.00750355783810508,-0.0138563822944677,-0.0191728376689088,-0.00308158727167684,0.00258075064404872,0.00354177556069457,0.00846818627780555,-0.00946023300048382,-0.0034907841597771,-0.00331121313906824
"946",0.0201318394048884,0.0291624068954848,0.0318932873085378,0.0181054698840277,-0.00600720621944961,0.000201476263923306,0.0130621973501777,0.0216829160069583,0.0196948300026172,0.0203488153415423
"947",-0.0000861320524448983,0.00566725345604291,0.0109671456446032,-0.000433657497820761,0.0125666697846607,0.0064516900127316,-0.00294716345628032,0.00757971935204638,0.00625996617070146,0.000406994849060593
"948",-0.00120654462926428,-0.00179300044983632,0.00394443816939516,-0.00889576528602809,-0.00833677189594673,0.0010019328214097,0.00221675120474818,0.000752327047804702,-0.0109248389488635,-0.0101708574073451
"949",0.00560879304637529,0.00487542265828766,0.00491186402117627,0.0120405503510903,-0.00439433576200654,0.000399802633873625,0.00129030970713817,0.0065142857945526,0.00989498388797205,0.0332921999423756
"950",0.00094380857135401,-0.00229846293578551,-0.00195502688515159,-0.000649429937955914,0.000192095753460908,0.000999601761628499,-0.00147235186085948,-0.00174268460827753,0.00478496871380951,-0.00477328649540332
"951",0.00308597958812706,0.000256118600312716,-0.00881505648417591,-0.00411238152708004,-0.00988122182023876,-0.00289649690341143,0.00866501737575964,0.00324199551534443,-0.00249441391987992,0.00479618003680238
"952",0.00777714052044232,0.0174000308104159,0.00296427051982184,0.0184743826171436,-0.00155016397625818,0,0.0098701470610314,0.00870016627028947,0.0159896929984249,0.00477332743478698
"953",-0.00390098792336069,0.00603617792656475,0.00689661525512442,-0.00170729169321193,-0.0149436157374295,-0.00571254454509251,-0.00307664675500208,0.00689979015786113,0.00507192484893348,-0.00158359108553852
"954",0.00204319207947967,-0.00249955187249984,-0.00782747270504625,-0.00128244591624904,-0.0122164554597286,-0.00433286764901519,-0.000545099356806467,-0.00587387951178875,-0.0079406827458256,-0.0111022708620921
"955",0.00492786058122885,0.00375949895570793,0.00690329766270792,0.00042810189831588,0.00807846379600563,0.00475645146863002,-0.00508586353343621,0.00787792755313577,0.00448837545944514,0.0100240858846563
"956",-0.0131042744027884,-0.0269664722141746,-0.00881505648417591,-0.03166475998575,0.00603509399816327,0.00342526489944972,0.00492955973820841,-0.0315095295327944,-0.0310544982950141,-0.0293767432883081
"957",0.00976581419328149,0.0197586736429429,0.00790513914633362,0.0159081353479531,0.00216393345198251,-0.000601512464566634,0.0199856543671548,0.0214377490308288,0.0092998692698496,0.0237218936144195
"958",0.00220590374049956,-0.000503092847206066,-0.0127452547605078,0,-0.0118737005258936,-0.00552604573409599,-0.00195963412020583,-0.00864190508365037,-0.0140877695810663,-0.0123852560833844
"959",0.00186253263692127,0.000755002168987495,0.00794439134026326,0.00108752014430946,0.00675221686305316,0.000303220068347931,0.00017848887955707,0.00498111715115601,0.00200814859034404,0.0084953217711945
"960",0.00295735658100105,0.00327055121771114,0.000985392655972417,0.0108626576419399,0.00286094424042815,-0.000303128153808396,0.0019630272965836,0.00272625715787966,0.00863339269662822,0.00521452919396115
"961",0.000168248739780053,-0.00802406314252424,-0.0098424261905129,-0.000859699928420832,-0.0154425418319589,-0.00666733835096633,-0.00587705045004405,0,0.000229262503816718,0.00518756107376728
"962",-0.00286410766471656,-0.00910020984359194,-0.00298203769927552,-0.0169930810302811,-0.00879122069394223,-0.00579679607842676,-0.0100325865331333,-0.00543717018439671,-0.0103912052876222,-0.00317590168457615
"963",0.000169263169910172,0.0104594090035539,0.00299095684534523,0.00634574018288392,0.00272155625513371,0.00583059484777526,-0.00615260280828789,0.00447292565411672,0.0132798096578193,0.0051772725314605
"964",0.000760068666843638,0.00025242294761485,-0.00397601117251867,0.00282687249908431,0.00934780770773003,0.00447469363701991,0.000728385421612909,-0.000742362986287715,0.010515010266877,-0.00237718728795866
"965",0.000337725423671387,-0.00630993256024492,-0.00998026666088914,0.0110582267151706,-0.00430591137326852,-0.00167444153798857,0.00727796864143637,0.0039614588380561,-0.00527821615435886,0.0063542032704953
"966",0.00793031314821158,0.0182878773641488,0.00705651542641195,0.0124380613175383,0.0131432493374704,0.00335440092405825,0.00559962007566273,0.0133169737508627,0.00432085361311185,0.0090765567807225
"967",0.00401776712846713,0.00698442899341267,0.00300316916057786,0.00614287858306262,-0.0203995036146616,0.00324271148939026,-0.00107785874515687,0.00219034841436572,-0.00694390493833852,0.00469301607448758
"968",0.0192582299717938,0.0240277100594695,0.0229540334125617,0.0227368151677687,0.00778366303509404,0.00807889652958393,0.0258948699086168,0.018212556831017,0.0338982424771019,0.0237446438397573
"969",0.00376235906604538,-0.0128205424629261,0.00878019571746247,-0.00185253314812683,-0.0171537320759683,-0.00420795525754913,0.00999137806612338,-0.00310037571347699,0.00257300597348387,0.00418253064980045
"970",-0.00187409340470412,-0.00833120754281169,0,-0.00412464881316366,0.00449081700896548,0.000301814720442994,-0.00485987968085999,-0.0095694503824415,0.0102653904434158,0.00265047491442716
"971",-0.00718433303527077,-0.0103778703630427,-0.00676965972900823,-0.0126321203261425,-0.0220476823156139,-0.00844750278528983,-0.0360999493075509,-0.0164250388800382,-0.0158949268100952,-0.00679756808052623
"972",0.00402933273781025,0.00124797968435497,0.0116846189963109,0.00734066906290942,0.00135039765054312,0.00375235203105428,0.0119412462346731,0.00171940446351626,0.01216910575025,0.0106463598290467
"973",-0.00376766111869875,-0.00997491842866027,-0.00577487536035493,-0.00978552280903389,-0.000518713568086415,-0.00111128299177943,-0.00804575919247141,-0.0132387008504484,0.00306032486664498,-0.00827682583247247
"974",-0.0118380652723009,-0.00554159794631948,-0.00774431972289813,-0.0241799597741282,-0.00539801576293353,-0.00829605033769421,-0.00937285285876899,-0.0134163154370347,-0.0288391826575858,-0.0417299075536764
"975",-0.00141438539838623,-0.00202610158148653,0,-0.000431068667820944,-0.0208748050865722,-0.0128527298475288,-0.0109171387749495,0,-0.00949961837834368,0.00158342810595902
"976",-0.0155792130638057,-0.0253809335346669,-0.017561312279526,-0.0262989670215612,0.0248374897292358,0.00744079358797367,-0.0314565469449588,-0.0198942585765239,-0.0109499850619239,-0.0296441914335533
"977",0.000507696594203466,0.00364583813557062,0.0148957960058975,0.00509234542138759,-0.00551324899373917,-0.00287218251759913,0.00873663617838449,0.00179892473229604,-0.00450481786283241,-0.00773932753243955
"978",0.0147182411012554,0.0238715384662407,0.0254401954088876,0.0237882138945151,0.00407965491913509,-0.00236619513436487,0.00696668792151511,0.0159011851807787,0.0131154389816137,0.0270935643193935
"979",0.00275094918575736,0.0038012487965442,0.000954364119759354,0.000645615940194411,0.00614500092846071,0.00206227291983474,0.00467424994257715,-0.00530143617106682,0.00083277313446195,-0.0143884167031987
"980",-0.000831296926097069,-0.0143903511693637,-0.00285960334517921,-0.00301013704415876,0.00424507883035652,0.00535031807852437,0.00204764110050903,-0.00380741773493931,0.00968229220156491,0.00324407562208728
"981",-0.0144769274580994,-0.0330428851458657,-0.0191207808841709,-0.03170142329773,0.00494908034502606,0.00204756245334781,-0.00705805920618996,-0.0236943009943082,0.00696739607334118,-0.00242518921933998
"982",0.0147739671404463,0.0105958694364474,0.017544086105463,0.0231620973082802,-0.0178504642727155,-0.0107252268523053,0.0192667336277941,0.0120043102265932,-0.00171126399192723,0.0186385273102563
"983",-0.011647269246593,-0.015202941909317,-0.0162835776479767,-0.0248145856734046,0.0138919232989454,0.00433669485303456,-0.00293602498452539,-0.0128934872421508,-0.00797430359084894,0.00477332743478698
"984",0.00303059570725739,-0.0167690734087479,0.00486870373652981,0.00781267939423858,0.00855038661362362,0.00215922877347996,-0.000552651041347496,0.00261259065774699,0.00300498833292018,0.00197938699468603
"985",-0.00562302027858963,-0.0151598121862326,-0.00484511431038304,-0.00819521302184234,0.0052099020121319,0.00174413519669492,-0.00386717681288762,-0.0122459513528781,0.0143060674970439,-0.00948249177806404
"986",0.021267964289535,0.0321606596085251,0.0204476308979122,0.0285842598025325,-0.0222288474702009,-0.0131506626140167,0.00758002869836405,0.0269059448148827,-0.000295325657883816,0.0295174429557872
"987",0.0128085653221444,0.0229029960198459,0.0095419806507453,0.0197568185073067,-0.00260714224473502,-0.00249687184715019,0.0135778503519741,0.0215771368625044,-0.00132964982531958,0.00852383101731813
"988",0.00269289050004895,0.0119758313138085,0.00567119776846603,0.00361932636858753,-0.00784273053942708,0.000104420826779528,0.00144833202277406,0.0057830751477761,0.0212278850864176,0.0126777038589156
"989",-0.00105824068927751,-0.0100335425796255,0.00469939803594466,-0.00169704532249904,0.0141223680220042,0.00625647327275103,0.000542048930187722,-0.00400003906707302,0.00753236725772033,-0.00113815050425914
"990",0.000570389431203244,0.00571760891581596,-0.0121608261519043,-0.00467467583516668,-0.0214071098042669,-0.0165805519618464,0.00325208673566757,0.000251086178580939,-0.018762137741628,-0.0068363323991949
"991",0.00366344914520478,0.00594283602454126,0.00284061922085765,-0.00640507632274445,-0.00966355895359594,-0.00853541378890565,-0.0149467108800054,0.00250957207103242,-0.0125275238095237,0.00764819747851098
"992",0.00389359685002644,0.00154154620563252,0.00188867906660661,-0.00343784793028856,0.00493199503865727,0.00212583849601833,-0.0107859886031154,-0.00150193007881827,0.00430300489740354,-0.00265651027620528
"993",0.00581775819525721,0.00461589769623605,-0.00282767802361938,0.00452798247467912,-0.0060815856391484,-0.00848473563748642,0.0103492358187363,0.00350948216758384,0.000295552939925781,-0.00152208837496137
"994",0.000642721329982887,0.0104678707549468,0.0132328598437195,0.00643909907506512,0.00375769549622906,0.00320957368598007,0.00256081990641666,0.00949301151251714,0.00472637900520279,0.00990851900668721
"995",0.000883197582557171,0.00151585563497991,0.00373132942354326,0.00149277844452422,-0.0145456351317322,-0.0105559466806551,-0.0102173816063814,0.00445436972989866,0.000955457531301773,-0.0026414734242225
"996",-0.00457211580817363,-0.0151362582137539,-0.00650563437048646,-0.0161842824191122,-0.0130238620205921,-0.00409458990043232,-0.0110596976048232,-0.0101012934783125,-0.010867940050489,-0.00264846928545504
"997",0.00580189741070791,0.00512292739496489,0.00561295005559659,0.00281413151252741,0.00692735111663789,0.00595126914450961,0.00260947946809931,0,-0.00660726815012469,-0.00341429533432092
"998",0.00107074095745974,-0.00713555034330482,-0.00279085150562774,0.00151122484362776,0.0182378060031674,0.0086042980815193,0.00780830752171413,-0.00971599636716725,0.00291457294543851,0.00761322130876096
"999",0.0024133173209917,0.00268690301074526,0.000932667267423692,-0.0045262168716701,-0.00107250503814871,-0.000106976044584206,0.011436843848448,0.00510755541755969,0.00678095395188438,0.00906686105773313
"1000",0.00634058321406084,0.00541078812778473,0.00591183452174238,0.0145972007018282,0.0069788445100305,0.00213372324214367,0.0109430236594454,0.00909300137775526,0.00155433349452783,0.00636464767940859
"1001",0.00311051484575953,0.00358799645364916,0.0037313036178479,0.00344071111781163,-0.00714367641188995,-0.00276677672981129,0.00696582620089536,0.00715627247160588,-0.00199529992634417,0.00520837720647793
"1002",-0.00143116160414669,0,-0.00092954876862561,-0.00107164780140123,-0.0020406109143426,-0.00352215835886782,-0.00307853146035586,0.00131551118326745,-0.00288781185736087,0.00370098782268258
"1003",0.000398189140016436,-0.0068948683030563,0.00279058686939515,-0.00321810110373988,0.0089317088270584,0.00385542704305619,0.0079924766203332,0.00630784523077144,0.0026733995938395,-0.0018437084596814
"1004",0.00143256460957297,-0.00128569851018201,0.00742145430056906,0.00086107785439693,-0.0195848924459169,-0.0105045506318467,0.00396499389939908,-0.000522415844552149,0.0162938596861544,0.0107130102608699
"1005",0.000715073399707888,0.00926870529859403,0.00920792458731179,0.0128025731809376,0.0169202321960986,0.0112432127358904,0.00448735878133766,0.00966813983650816,0.00357095173028021,0.00036549207135006
"1006",-0.00158823415747222,-0.00459174149799735,-0.00821164668886076,0.00509894566422031,-0.000751975989216613,-0.00203125686285754,0.00125090729466715,0.000776631768113711,-0.00493797084768133,-0.0120569444895691
"1007",0.000238669908035005,0.00666332405339976,0.00367981432649755,0.00697489926447781,0.0110647485589623,0.00503465147949256,-0.00124934448054281,0.00672314287965148,0.0123330804373718,0.0188608017722003
"1008",0.0103380446955743,0.00814673777567987,0.00916602216017526,0.00965606091317772,-0.00754392127310399,-0.00309116886476191,0.0155469206556982,0.00899040514377902,-0.00519031859003516,0.00435584443840731
"1009",-0.000551175467547571,-0.0020201670861304,0.000908415289868403,0.0045734936944748,0.00117781727021438,0.00235249170790408,-0.0177720477502258,-0.0050914499125877,-0.0235507246376812,-0.0133719597444494
"1010",0.00519787716744191,-0.0063261143630764,-0.00725950371814221,-0.00248309929310664,-0.0220274403821472,-0.0107731697695931,0.00411998767261634,-0.00230295078955145,-0.00282007421150288,0.0106226410499182
"1011",-0.00195857078633244,-0.0114590095260151,0,-0.0105809006028412,0.0043730928414778,0.00517574868289294,-0.00535198176927132,-0.0143625524877665,-0.00401870224077916,-0.013410585848192
"1012",-0.00196271125442005,-0.00540922239964636,0.00365594663037716,-0.00922609093549831,0.00533415774826418,0.00665062442032238,-0.000358873974525165,-0.00312286316171351,-0.00186804151732733,-0.00367371914114689
"1013",-0.00125849107892839,-0.00492153314507571,0,-0.0103707716924343,0.00541492250535147,0.00341024690514069,-0.000358925116266007,-0.00313238946801975,0.00404246887194981,0.0117994381284996
"1014",0.00354372716893847,0.00702753072077433,0.0072861658791219,0.0106926908283165,-0.00560081487773278,-0.00392971887012605,-0.00179524404116493,0.00418980013778869,0.00589031486319391,0.0112973335278741
"1015",0.0090248772889252,0.0294651507302361,0.00904141654112478,0.0201019208133202,-0.00779807187862513,-0.00287871389310823,0.00449592230423335,0.0151237539962854,0.00407681405153615,0.0064864718915163
"1016",-0.00163364202868166,0.00477055266571735,-0.000896021806504832,-0.00871203120924358,0.00895144931347658,0.00673676272402024,0.00286420159605361,0.00154135655785259,-0.0104090058108441,-0.00143220592840976
"1017",0.00724495937320158,0.00924509054665124,0,0.00292967885378626,-0.00638354671339481,-0.00276203555490184,0.00678308941221006,0.00641201506773115,-0.0101454753417649,0.004661289919627
"1018",0.00170144005020001,0.0099035362364297,0.00269055496581383,-0.00146061192822022,-0.00468197871733955,-0.00244962832833673,0.00939746462790758,0,0.00557684067259268,-0.00107079602915094
"1019",-0.00980539820485049,-0.00833554384702839,-0.00178891640629009,-0.00773095965535098,0.00721995774111139,0.00256304435124943,-0.0119448030688217,-0.00535179367816507,0.00217348433796283,-0.00107179677897651
"1020",-0.00132571295129147,-0.00642769429979939,-0.00896040181593116,-0.0109496521468759,-0.0137933657765609,-0.00777445936585397,-0.00213292445994751,-0.0102485000774871,-0.0188453782617007,-0.0100142801895847
"1021",0.00226410443659963,0.0126897314876897,-0.00994564560387035,-0.010432021086229,0.00792915248535953,0.00332749400883015,0.00391929411769554,-0.00025901494103675,-0.00129571649304228,0.0101155804464559
"1022",0.00568703697922879,0.0100738088757368,0.00639273300927123,0.00774525214095712,0.00043690188937151,0.000106440522863904,0.00496881876875599,0.00699127115304843,-0.00511331759988787,-0.00858361088916537
"1023",0.00054228154242919,-0.0026757263647913,0.00907402076902541,-0.00597782650955969,0.00950251822772041,0.00502770996211477,0.0105948177428272,0.00539953815350613,-0.00199443846276126,-0.0126262752838782
"1024",0.00387067761131599,0.00536574492754127,-0.00179838455728676,0.00880571380502815,-0.0151469152505789,-0.0060660536881435,0.00279599134142017,0.00332504470318318,0.00814756303700692,0.0222871715082313
"1025",0.0024680238520558,0.00557987424338546,0.000900759501514914,-0.00340623702021481,0.00450429834735,0.00374775962694196,0.0139398964364383,-0.0025488231842582,-0.0246264402370709,-0.00857762194444589
"1026",-0.0174631777978554,-0.0243667804703982,-0.0171014806650615,-0.0316173056905438,0.00524891413378414,0.00458680712352888,-0.0156383221823908,-0.0171222892638666,0.0183694129602125,0.0126171730460689
"1027",0.00751653305653521,0.01409515269859,0.00091560710116223,0.010588931573438,-0.00761456207029443,-0.00392861887656959,0.0118713115857831,0.00832013015739386,-0.00314709858111084,0.0156639803234693
"1028",0.0160084467435508,0.0246282109307985,0.0201280655902352,0.0242306557695111,-0.00495094519773598,-0.00464961220973392,0.00465837542627723,0.0180506941413208,0.00716106903677027,0.00736068056253858
"1029",-0.00191171165705717,-0.00333180034062808,0.00986555212365992,-0.00745958243701084,0.00022106144483125,-0.00236211455341073,0.000171423057506725,-0.003039559072891,-0.00267588678877939,0.00974249329415966
"1030",0.00222228824152371,-0.00501456719282767,0.00799265529798521,-0.00128836316000813,-0.00828953934298171,-0.00570447943103936,0.00257593593623562,0.0015241009859841,0.0134151018799946,-0.00654715488960811
"1031",0.00282906433470598,-0.00287955998669798,0,-0.000215101447783805,-0.0101432544792968,-0.00617032274612295,-0.00907718581581873,-0.00608820682801547,-0.00408466726364609,-0.0055498412586894
"1032",0.00625234004407482,0.00601671907424972,-0.000880738512264112,0.0012904884277849,0.005179383714913,-0.000436002101953603,0.0112342094699627,0.0028075383156243,0.000151822872495266,-0.00279037104622348
"1033",0.00454682568886211,0.00717692640382794,0.00617287761848839,0.00042966139359768,-0.00918528534161367,-0.00686450886556322,0.00256365360958921,0.000763700163978642,0.0110875309660747,0.00664576963206298
"1034",-0.00226319185288482,0.00190045929089888,-0.00701167861682195,-0.0229715169736184,0.00870560168395595,0.00570526364629997,0.00238648874314129,-0.0094097953612462,-0.000525702272237361,0.00486435090443704
"1035",0.000378164955475935,-0.0101945697873856,-0.000882370721157488,-0.00944821019128828,-0.0115446110745699,-0.00327280867551094,0.003231282782028,-0.00744572544016742,-0.00165327262664072,-0.00587820501003333
"1036",0.00597036284274655,-0.000478857533316668,0.000883149986848242,0.0122006061637281,0.0144004277687413,0.00459668076781061,0.00627246249185465,0.000258983426713044,-0.00398945409155649,-0.00347824910264893
"1037",0.00240389313532163,0.000239415272906163,0.00882644797511101,-0.0050406896175107,0.000670234107593037,0.000327306183178333,-0.000168524496668376,0.00206849318549729,0.00476110917980832,0.00488653099623337
"1038",-0.00314781887931925,-0.00167704381183242,-0.00699951200408433,0.00198251103718183,0.00446918847067979,0.00228757577827676,-0.00336981778558254,-0.00567759694425463,0.00767208742396597,-0.0128516878535987
"1039",0.00631531603675639,0.0112793464943308,0.014097210632501,0.00835336223772409,-0.00322480911924072,-0.00141356252004377,0.00287408741758455,0.012457931007277,0.000970403814507748,0.00738913410732644
"1040",0.00298862369707065,0.0042715131633444,0.00868782759616549,0.00348802842487683,0.0015614564393267,0.00370074120730268,0.0013484238064394,0.00845961363396475,0.00700959700180781,0.00314354882990564
"1041",0.00208549750835285,0.00472591073522022,-0.000861014804973137,0.00608312744562833,-0.00311902508655482,-0.000217008293725174,0.00387214192655527,0.00279586935428844,0.00274001050933093,-0.0010444823480118
"1042",-0.0200698441114835,-0.0275167478498235,-0.0275862938066121,-0.0319584584498193,0.0149737363265112,0.00965214775043166,-0.00905572959807421,-0.0240810915513759,0.00649870005173336,-0.0013942307795789
"1043",-0.00614417053961525,-0.00096701191377957,0.00177287521694769,0.000892126396377479,0.00363355860565995,-0.00247115758971683,-0.00795430283516696,0.00545440514303119,0.0089515156112745,0.0223385505785685
"1044",-0.000686961963731525,0.00145209996493034,-0.00265463246418185,0.0024515526114981,0.00636197147135897,0.00258482753230682,-0.00545867113071752,0.000258479712790916,-0.00749035733729753,-0.00887669868527741
"1045",0.010692625679368,0.00991040204102922,0.0133096871942386,0.0120054227238808,0.00588614304219526,0.00322154224393545,0.0178387278608065,0.0178202123740492,0.00659443893887568,0.0220461048357377
"1046",0.00619673492975847,0.0117285493906696,0.00963212236685607,0.00593128438425738,0.00130057091698221,-0.000428521143521432,0.0208969328925945,0.0134486134562937,0.00203813502554451,0.00168514618857385
"1047",-0.0166729202760706,-0.0160870964703399,-0.00173453640393462,-0.0102640457532319,0.00289896051350524,0.00113825404572321,-0.0269068289614625,-0.0160243037884985,0.0172162932669973,0.0151413553204189
"1048",0.002138379747747,0.00673214232079133,-0.00868803121135853,0.0136800978156961,-0.0153730561914291,-0.00525413775391781,-0.00797292434633945,0.0050890667957626,-0.00078555310137518,0.00397754323492205
"1049",0.0172242521657666,0.0128971774361637,0.00964035845536149,0.0198087240574694,-0.00978562049650622,-0.00679087452679095,0.0143639687020836,0.00860773325157527,-0.0130789167106762,-0.000330205386527171
"1050",-0.00749236571233203,-0.00848860727350542,-0.00694424577404229,0.00106709633836433,0.00832795800221775,0.0071628799604242,-0.00859767379131771,0.000501844330330847,0.00912455671300028,0.00495373116318754
"1051",-0.0078503499690773,-0.00808571223284227,-0.0192306441473103,-0.0140724086622237,-0.00638700205254872,-0.00247816928386158,-0.00646129511816662,-0.00777704814619273,0.00265514879131024,-0.00460062643848858
"1052",0.00874971397410174,-0.000239369800400513,0.00445625452008636,0.0134082383574889,-0.00609596052652672,-0.0023766657497164,0.0124933799699629,0.00227550031956048,-0.00257658171645725,-0.00858377702770841
"1053",-0.00143331138020852,0.000719275608060732,0,0.00192055854252349,0.00970139811252846,0.00584796154130984,0.000507477962609304,0.00327962408650739,0.000358804532442303,0.00399601803386762
"1054",-0.0185059527094718,-0.0230051796068057,-0.024845056157371,-0.0296059450829801,0.0167864633371213,0.00850379983244798,-0.015543416931374,-0.0226302798447117,-0.0117638616522814,-0.0162520558719252
"1055",0.00692621124085968,0.00392468226466258,-0.0163783587190829,0.0103161059783217,-0.00564821094213452,-0.0023481195171603,0.0113266406820454,0.00102915720688146,0.00326629155066294,-0.00573161612253437
"1056",-0.00603746999353094,-0.00464240787358849,-0.0703053019759884,0.00586567572572561,-0.00043629500117881,0.00224702417286382,-0.00678784110282293,-0.0187614200497178,0.00463029948900107,0.00271274688097622
"1057",-0.0114573532887132,-0.0252822332494375,-0.00198985426177256,-0.0166307150989816,0.014970625355204,0.0036302567250095,-0.00802994066034779,-0.0275013353276056,-0.01865185785214,-0.0365235273160286
"1058",-0.0185128634813625,-0.0307226365067208,-0.0368893227437794,-0.0204258328990863,0.0113053329166226,0.00850898731964844,-0.0130900148893108,-0.0250468003918185,-0.000220143825636065,0.00596703307699742
"1059",0.0132351622562836,0.0350741291112933,0.045548567786305,0.0123318024721024,-0.00766601213117524,-0.00305853117177879,0.0083770956246525,0.0256902591856558,0.00535816187029647,0.0310536687711132
"1060",0.00363698793585909,0.0107930451996492,0.0267327704200091,0.00177193496970807,0.00268248730869591,-0.000635045856788086,0.00882645171784913,0.0237395478242703,0.0102211724449064,0.00575298742614816
"1061",0.0154982287640741,0.024584226022794,0.0289296662227572,0.0192347742511221,-0.00588474466533007,-0.00518699439496528,0.0109796921700673,0.0237966894822226,0.00556481916473284,0.00471070698178733
"1062",-0.00346877024703773,-0.00266586890386011,-0.00374898084784669,0.00303699899383947,0.00333622550768853,0.000531718216735033,-0.008993616987509,-0.00723131869704363,-0.000646801787025919,0.00736764965761338
"1063",0.0028618261808071,0.000728889245399378,-0.00564426084688308,0.0131920943474206,-0.00128785989269631,-0.00127594840967937,-0.00753430010040435,0.00884510428749374,0.00927718786169329,0.00199472211951734
"1064",0.0095635009095314,0.0150557056431924,0.0018920443563244,0.0115261254947634,-0.00751774851613973,-0.00511171420086265,0.00465837542627723,0.0105723659306842,-0.00798058309763683,0.0033178730098975
"1065",0.00305577966673143,-0.00885165881892147,-0.0245513715393736,-0.00105524936777179,-0.00248996505457788,-0.00267645065042843,0.00507542131194616,-0.0109719785829773,0.000287271941622924,0.00264546644963271
"1066",-0.00243715035051095,0.000724189307791834,-0.00193600280915662,-0.00506957830098531,0.0014106581030735,0.000322764551589971,0,-0.00438622787093901,-0.00517019981222888,-0.0135224126400227
"1067",0.00671857929159114,0.00410011374509089,-0.00194024122934755,0.0114647638984016,-0.00769203897508963,-0.0028984954717739,0.00448144765260006,0.00103672458543591,-0.00238188260916128,0.00568367458562014
"1068",0.0069012807901816,0.0100890117148746,0.015549314655958,0.0128043942121585,0.00797014709604738,0.00344440878613983,0.0116675169993496,0.0111310746356692,0.00332820328993977,-0.00132973490910149
"1069",-0.00135581598461321,-0.00546967260748654,-0.0124401159784582,0.00870491303306609,-0.00205788793589612,-0.00257396383808772,0.00746280645884956,-0.000767916237635946,0.00858154624044927,0.01564586580112
"1070",0.00422362337899118,0.0119561965383157,-0.0019379922529702,0.0160262269054654,0.00486168039562362,0.00213401695462379,0.00235677898729869,0.00922345448422179,-0.00471903328529233,0.006882928416728
"1071",0.00082607046298655,0.00543449079242553,-0.0135925150537165,0.00849347039813275,0.00108404326681022,0.00225889781009392,-0.000839547490751658,-0.000253855208783182,0.00459769406460553,0.00911459275608784
"1072",-0.000149968713895166,0.00258520479306767,-0.0196848932712549,-0.00200495145387536,-0.0040091974887837,-0.00504396535602381,0.0016810590395353,0.000508129008902625,0.0158038262529698,0.00096772869811601
"1073",0.00315210412433609,0.0114863576909714,-0.00903619675943435,0.0054246953714705,-0.0150129824576468,-0.00431454062059744,-0.00134272472270291,0.00736009601031573,0.00232313969046527,0.00290047881931033
"1074",-0.00254377454525267,-0.00370771440844753,-0.00810537416792678,-0.000999267245106794,-0.00198750940790748,0.000108377830452033,-0.0104184489143496,-0.0136053474903871,0.000912979318971052,0.00192792795831886
"1075",-0.00345043465886086,0.00790838173976427,0.0194076552895202,0.00100026677893528,-0.0053129459852127,-0.0029251024591177,-0.00747148224443273,0.0107279445331034,0.00806967258682434,0.0237332348437118
"1076",-0.00301056284931278,-0.00138459017834569,-0.0070142770343542,-0.0117906139334264,0.000890742672970735,0.00130321470955042,-0.00102646462825551,-0.00732855978253588,-0.0071001320590246,-0.0184837784171399
"1077",-0.00747394927716283,-0.00970640404259893,0.00201829051576685,-0.0188070075864305,0.0107827025996738,0.00564294619652084,-0.00205503868102708,-0.00789200359362952,-0.00722096191265387,-0.020427623687187
"1078",-0.0000761392852290932,0.00093325424913937,0.00402824393664347,0.00824416732865041,0.00626847650944096,0.00388433336312022,-0.00120144988245163,0.0030789672360485,0.00204782852872087,0.00782006312591998
"1079",0.000760887064799709,0.00349728231863922,0.00702098974608467,0.00306643508973092,-0.000765006567203019,-0.00333221572525877,0.0135740693696877,0.00818629394625892,0.0134602119856329,0.00258645032519977
"1080",0.00364835255074336,-0.00232327167515001,-0.000995859697986878,0.00122272376739896,0.0135624460482608,0.0073332774066317,0.0110187346844615,0.00304521262464008,0.00862252289301879,0.00515972166490997
"1081",-0.0112086978273926,-0.0251511280685617,-0.00299111221216952,-0.0250357784542473,0.00226532240134936,0.00246170489540876,-0.00989292590049673,-0.0146724822925601,0.00606680442467833,-0.00609568631687829
"1082",0.00574472988834351,0.00859975368568855,0.00300008580545974,0.0144048892580084,0.00430703595049109,0.001281937084743,0.0077900860274922,0.0077021867964806,0,0.000322850943261122
"1083",0.0136316661412894,0.0272382448983175,0.014955298193229,0.0236675296594642,-0.00643206198431878,-0.0039462947763077,0.0115947684508619,0.0168149891577272,0.0039060304758598,0.0158115350310737
"1084",0.00510902697335314,0.00691752197436357,0.00392908713551798,0.0088459443093043,-0.000863415349978913,0.000750189933567347,0.00714287496902699,0.0107743657900208,0.00163825938566542,0.00730619171549063
"1085",-0.00104673567582458,0.00160301805106555,-0.000978520616824685,-0.00817024622838003,0.00377963765654732,0.00353043013908771,0.00494771531365457,0,0.000885852498096806,-0.00283811777633758
"1086",0.0086052595759345,0.00983039441563438,0.000979479057275912,0.00863939943280423,0.00968319110621185,0.00426460283583951,0.00935517943964181,0.00793254677111821,-0.00333621581453702,-0.000316316289468599
"1087",0.00652879742931312,0.0178856144767259,0.00195686924654792,-0.0017926043135541,-0.0102295953941716,-0.00286663068579984,0.00455288670326759,0.0108217511390414,0.0192648715922641,0.0060107715714699
"1088",0.00324288853838484,0.0040036236265375,0.0263670552134689,-0.00818205148877527,0.00764356605857763,0.00383325643186061,0.0111688313733642,0.00389289038100293,0.00415556308623799,-0.00723270247891861
"1089",0.00235122957599998,0.00443052431046254,0.00190298569346226,0.00603614753645076,0.00309796371992999,0.0020153601115096,-0.00480241952653049,0.00484711482661515,0.0170203436180589,0.0104529163490235
"1090",-0.00153917433654216,-0.00220556442112985,0.00284897336387258,0.000199988655960492,0.00160472175734938,-0.00030794984918614,-0.000160668247342066,0.00144720263305254,-0.0128633659140043,-0.010031372377705
"1091",-0.0035971720308422,-0.00773664238146277,0,-0.0221955848739055,0.00566019093036818,0.0026542538510046,-0.00675695412719601,-0.00939273260417717,-0.00352369513932049,-0.0104496070956075
"1092",-0.00663103615874683,-0.00757389634790584,-0.00189364243259305,-0.0165643359418466,0.00446012905198012,0.00254081191524569,-0.00550697766343977,-0.0111845142542076,-0.0143448687501713,-0.0160000118565692
"1093",-0.00904787797318318,-0.0255893109634149,-0.00759024679954845,-0.00956541954799006,0.00951450197362336,0.00496338488533365,-0.00146589610333203,-0.0118023932473813,-0.0288363576480433,-0.0669918253132131
"1094",0.00441567350401195,-0.00483745834928639,0.00573632948458913,0.0130167336211282,-0.00439838150562033,0.000525409701298996,-0.00538204957850319,0.00870888525660507,0.0127552937007369,-0.00313697441194594
"1095",0.00387483448361792,0.00555527399482791,0.00380190654496659,0.00186543529461147,-0.00105185504556482,0.00147062917293805,0.0039355327703583,0.00419340008294422,0.0143152233795893,0.036713179193959
"1096",0.00853599224202384,0.0112802968686174,0.00473485510500593,0.0117914217818667,-0.00715992203181959,-0.0048241841776141,0.0138842887821562,0.00245668074174632,0.00352821944876425,0.00910628911108069
"1097",-0.0105247466938982,-0.0168451606122791,-0.0169649244377231,-0.0220812345144626,0.00572659848441415,0.00358305450443064,-0.0111163711003996,-0.0161726964957647,-0.00919540943321462,-0.0320855705109503
"1098",0.00476059153195818,0.00324145098463169,0.00287628801696926,0.00292704777478092,-0.00632684743282352,-0.00220557430127954,-0.000162736122689244,0.00547889504965404,0.000341224255415495,0.00103589746505772
"1099",-0.00769898530669189,-0.0159242532219956,-0.0210325639532303,-0.0218887502067545,0.00902038677823791,0.00389461432467719,-0.00912515132073199,-0.0118895785705984,-0.00654881660546602,0.00172481566061466
"1100",-0.00634154183046887,-0.000468925322591685,-0.00585911355599633,-0.00149184287197757,0.00557425081113361,0.0024108972444763,0.00230203780758553,-0.00200538579757248,-0.00178541503174445,-0.0130854680616797
"1101",-0.000150193465877302,0.00187695783833397,0.000981933652456357,0.0032014996591252,0.0102500719189857,0.00292816895143355,-0.00147653115748114,0.00728429474892445,-0.00433370036230651,0.00244246696417449
"1102",0.00893576894047121,0.00702578136983179,0.00785083937050923,0.0161703751143725,-0.0132520073591108,-0.00573520877452349,0.0111732568591032,0.00798014609128805,0.00594169524866328,0.02018793134022
"1103",0.00238185342820629,0.00837210453883608,-0.0146055822734668,-0.00649101350976133,-0.000419644959684051,0.00104846104451495,0.00194984887869043,0.0056905308202817,0.000343324161676151,-0.00784711418311368
"1104",-0.00794450031390592,-0.0161440499873133,-0.010869539101471,-0.00800821190282408,0.000524272634021772,0.0024099491445535,-0.010217353958728,-0.00787225088189947,0.0126331004174296,0.00928471077985238
"1105",-0.0116014047449767,-0.0241444478304108,-0.0149850637224885,-0.0208200548972479,0.00482572205268017,0.00135874605068542,-0.0104864719049746,-0.017604998528169,0.00230522061478,-0.0160136901516122
"1106",-0.000832879656341712,0.00312302417510124,0.0121705563096728,0.00998038925000855,0.00375887528924501,0.00104427871227664,0.00298046932873097,0.00555296999740262,0.00514099972751136,0.0135042207483271
"1107",0.00333459033911487,0.00933903904527145,0.00200392819004858,0.00214826517106603,-0.00468013682271906,0.000102981623234522,0.00412744041904256,0.00301222203538121,-0.0000672589021404324,0.0181072403749749
"1108",0.00460780727545851,0.00972719537604982,0.00899984728444481,0.0128620923423877,0.00856966769284706,0.00552626146253066,0.0129893267778789,0.00725731802098784,-0.00242294383600838,0.00369129388523048
"1109",0.00383432206929646,0.00798863086636947,0,0.0105817993729582,-0.000414625840659877,-0.000103362972594168,0.00178531901699763,0.0111799267654531,0.00998513014448021,0.00568367458562014
"1110",0.010411276929696,0.02191159075676,0.0178394643605282,0.0163350297546934,0.00228039964248183,0.00155467312568924,0.0174985981314044,0.0122852603942194,-0.000400788251184836,0.00565158721344039
"1111",-0.022460983683953,-0.0278285484745997,-0.0126580115638507,-0.0179271318071036,0.0135147942804401,0.00824140404825524,-0.0281849951051593,-0.0177186434689909,0.00180436381852678,-0.0125619145801649
"1112",-0.0010616202530539,0.00821227109042777,0.000986125113052738,0.0094418888136325,-0.0190496316034049,-0.00597094378555307,-0.00573478346178735,0.00716558060168815,-0.00273500092762313,0.00870430105841091
"1113",-0.00994462606954594,0.00744686397335936,-0.00886716193440029,-0.00498872120445615,0.00574243604920288,0.00393610274676681,0.0036255987988052,0.00147213655426914,0.00481606020066883,0.00398275562528294
"1114",-0.0105813244713194,-0.0157081155306562,-0.0099401680201644,-0.0160850695468959,-0.00757812388200296,-0.000619484051193164,-0.0142857515421136,-0.0100439674336067,0.00173076153820562,-0.0115702605873167
"1115",-0.000619492629924556,0.00938749510420567,0.00803201476098403,0.00785552178084092,0.00460213119269293,0.00185849234422575,0.0119939698002816,0.00296937014365106,-0.00039871080273024,0.00936459327804839
"1116",-0.00418761546846391,-0.01697297977048,-0.000995859697986878,-0.00716242914296328,0.00780928909650025,0.00216323244668648,-0.00477370674198496,-0.00764848430750731,-0.00405531184756425,0.00828362085452339
"1117",0.0076311827909481,0.0130088868120561,0.00697898922493945,0.00785091495942325,-0.00402908454936601,-0.00400960350004209,-0.0092623104222006,0.00372896332364214,0.00500634143256584,0.00558665132076031
"1118",-0.0139105260734997,-0.02638330080095,-0.00990100244771031,-0.0216841989682147,0.00767606832655776,0.00320040327371562,-0.0237061055949044,-0.0173391840402503,-0.00876722248628092,-0.010457541356911
"1119",0.000783609357947412,0.00263773946680268,0,-0.00172178803151724,-0.0050440809659591,-0.00216137321587917,0.00188087404600812,0.00252079831140528,-0.00984991256198364,-0.00660506552415063
"1120",0.0126862958049045,0.0141113646623352,0.0199999373084043,0.015089535775034,-0.0151055547841318,-0.00793989759855351,0.0157023222146557,0.0145838590230649,0.0060905053504634,0.00698149320234909
"1121",-0.0177855163069366,-0.0360849240733185,-0.0196077828800465,-0.0214480968473345,0.0181735093592821,0.010809415108596,-0.016467752196763,-0.0195788372518215,0.00302681782507319,-0.0267415394978376
"1122",0.00220459929511052,-0.000489462629133852,-0.00299999792004524,-0.00759566994904926,0.00454004609754488,0.00277633362305041,0.00700479545289312,0.000505569836483311,-0.00100586108522871,-0.00407053551353975
"1123",0.00298404119194662,0.0124848390198162,0.00300902498875288,0.00131200159780565,-0.00472478644515373,-0.000717672812352355,0.00848307566466611,0.00319184270358042,0.00651138479887625,-0.00442780233597684
"1124",0.00511631769002951,-0.00362671899217348,0.000999960246497622,-0.00152855067242863,0.00123878353827989,-0.00153908356827959,0.0105992495415883,-0.00254516922252035,0.000600220080029246,-0.00547389412708488
"1125",0.0137037433397684,0.0232684010783255,0.0169833082968665,0.0183725772869932,-0.00443227626554576,-0.00133640167385651,0.00882277958276578,0.0130135503897404,0.00486566689905787,0.000688055927610343
"1126",-0.0060254100101963,-0.0126058198746577,-0.0011892154090547,-0.00995695305239896,0.000620976877493185,-0.000411014630463113,-0.00214501994214267,-0.00881617528579737,0.00152566998957515,0.00446882846379237
"1127",-0.00287570150195671,-0.0122759696253172,-0.00198392456113827,-0.0013144449817748,0.00765671508903298,0.00525081905892022,-0.0183561355935909,-0.00304963630487953,-0.0175508902062754,-0.021218265704642
"1128",-0.0116133989333419,-0.0156601346673629,0.00596360502589843,-0.00175531090340786,-0.00421034696944711,0.00419938661413433,-0.00108795969099107,-0.00994115338671475,-0.0140218488343495,-0.0118882007975992
"1129",0.00891103579307795,0.0111111727823991,-0.00494025244363139,0.0116484904842771,-0.0137141728552466,-0.00387600499512131,0.00527576980518485,0.00437688408350412,-0.00362367713741552,-0.000353779382827213
"1130",0.0130529866317985,0.0119879173900805,0.0119162615173323,0.0136866690195445,-0.00804964632285177,-0.00921459119221879,0.00829529290729991,0.0125606529436333,0.00349968444382576,0.0176990911858448
"1131",0.00856424757398155,0.0194966310149394,0.0157019230158115,0.00921558636960262,-0.00664000757177574,-0.00599311703452943,0.0110811845050964,0.0091140041476836,0.00642770765769596,0.0180869597716493
"1132",0.00956220381348372,0.018639760005303,0.00772935354028315,0.0108303299660448,-0.00159196646582038,-0.00343181163535244,0.00132826467983582,0.013045589129884,-0.00801734648811947,-0.0105910798016576
"1133",0.0147760955053509,0.00879252192743962,0.00862909199816841,0.0117647716902394,-0.00159936996052579,-0.00249873978078829,0.0179106791864709,0.00841996180313953,-0.00732881506849314,0.0013812676985363
"1134",-0.000820979380500964,-0.00777380996666466,0.00190125037510169,-0.00041533178636588,0.00224304962666544,0.00628994563177399,0.00619085213946202,-0.00736760386393709,0.0186297669937789,0.0134482335920072
"1135",0.00119540158934939,-0.0104462459933325,0.00569223859540835,-0.00664728322892527,0.00511525442161243,0.00177137736860389,0.0061526235519942,-0.00395817079656979,0.00867031739245672,-0.000340247139329009
"1136",0.010375562670625,0.00791717178825757,0.00660390967036473,0.0138018920153444,-0.00296937854231871,-0.0038481413424053,0.0125525596077154,0.00596153115956533,0.00161164457426244,0.0211027479228436
"1137",-0.0070925934663878,-0.0147580517199202,-0.00843499790051838,-0.0113452378283093,0.014143699647861,0.0106478877403415,-0.00349665951077716,-0.0069137894314838,0.00737516623701651,-0.000999986380040063
"1138",-0.0180801608814123,-0.0374487655479803,-0.0122870035093764,-0.0279572034637078,0.0149941377542921,0.00764431849917058,-0.0188198299504913,-0.0236200602803999,0.00891844259567387,-0.00767430506191968
"1139",-0.00431912452023697,-0.00803216346336522,0.00287058971052123,-0.0100881402490551,0.00340915542023223,0.00143499487768461,0.00341383528330619,-0.00127339704356388,0.0077842076069452,0.00874238413852768
"1140",0.00334846077237416,0.0156880941200899,0.01908404784121,0.0162619954882388,0.00277945265305601,0.00163752541248474,-0.00842388246490688,0.0104540098928709,0.00896769630247563,0.0136667549848453
"1141",-0.00690207796666997,-0.0072248573893775,-0.00936348317429914,-0.0106677455654578,-0.0142707903954762,-0.00572240832624249,-0.0111093809461551,-0.00782215459406888,0.00259500455816153,-0.00559029126745914
"1142",0.00580471359952139,0.00150588921267469,0.00756149053479627,0.00625403704731653,0.00166603925343733,0.00411108532831839,0.0109038905153134,0.00508641287546885,0.0042707650439715,0.00892861944212275
"1143",-0.00820112931979777,-0.0175393841025397,-0.0121949834064761,-0.0115732025722068,-0.00967049669068953,-0.000613992590364987,-0.00898846082332183,-0.0129048834607496,0.00882738419125095,-0.00557203579296839
"1144",0.0162314031765753,0.0132618015869919,0.012345537025648,0.014527554242403,0.0207898294789466,0.00378972461694804,0.0173151940627394,0.0115353854721298,-0.0121990350297424,0.00692156308141456
"1145",-0.000602559823581816,0.0135918937978319,0.0103190291068784,0.00299184767450367,-0.0118284203667081,-0.00489775474183352,0.0074567246062327,0.00608218849594477,0.00879348225026555,0.00327327776015629
"1146",0.0138710140612948,0.0273155899514996,0.00835657067316631,0.0159814218453218,-0.0077031881464672,-0.00553749895064459,0.00643608823434749,0.0118387223725065,-0.00762723990187819,-0.00489389755420977
"1147",0.000669087337975105,0.000483572696178047,0.00184175379481477,-0.000629102976362428,0.0075528574640118,0.0038149404909269,0.00511564469420911,-0.000995781077172797,0.00833167334067442,0.00819671052420667
"1148",-0.005572712331815,-0.00579851874039294,-0.0036764156322272,-0.00209880845290611,-0.0109318173713875,-0.0031847587217908,-0.0112929217054453,-0.00647882778197728,0.00781450832098751,-0.00487801563658707
"1149",-0.00373632233338528,0.00680392232918337,0.00184483002053026,0.00336497140388192,0.00684197782234053,0.00422606126808267,0,0.00476512532346729,0.00273298595990812,0.00784313079179988
"1150",-0.0204754511678943,-0.0263091163593653,-0.0165745540176513,-0.0176064693143101,0.000104727006642102,-0.00164201083716131,-0.0268660897966602,-0.0154762677235921,-0.00367625014448247,-0.00680941221417808
"1151",-0.00290968613717379,-0.00421442595546195,-0.00187279452889799,0.000853604140682362,0.00376338713264923,0.00195255875319877,-0.00148810831883361,0,0.000827056418003069,-0.00326472866915961
"1152",-0.00683451502502896,-0.00199116249027154,0.00469053960044508,0.00426336518876136,0.0197877538348754,0.0121051615401453,0.000496931865941352,0.000253287203852759,0.00616568749580604,-0.00818865621833109
"1153",-0.00425274111857565,-0.0164630303444858,-0.00933714672536745,-0.000848944324963519,0.010092080795155,0.00363771567874394,-0.0132386697184516,-0.00481606154460923,-0.00360093515197779,0
"1154",-0.0255474873293534,-0.0304339027449902,-0.0084823975285534,-0.030805277263064,0.0300262979862891,0.00921259896920446,-0.0293479075550435,-0.019103722698692,0.0240933488201032,0
"1155",0.00541887131422203,0.00706273137589974,0.00190125037510169,-0.00350724926826229,0.00196990028097899,0.000802312127015758,-0.00621947937117417,0.0111663096772299,-0.000185729316846794,-0.014861261469488
"1156",-0.0468417391644634,-0.0727272059987167,-0.0607212529344988,-0.0571931435728162,0.0355810833385812,0.0132301637912042,-0.0483307592317427,-0.0606063053058453,-0.0052635207980829,-0.0378813261809202
"1157",-0.00149660764878279,0.0240896539008755,0.00909105310032543,-0.00653282014888057,-0.0288532683891874,-0.0115742485388126,-0.0206429839728938,-0.00328048029366645,0.00690986682588313,0.00418112739105347
"1158",-0.0651236509406113,-0.0820570044026349,-0.0480482015217951,-0.0833726497087643,0.0315679199801711,0.0159132699835103,-0.0850592071041384,-0.0811850013429679,0.0331993508500772,-0.0371269529125423
"1159",0.046499632136165,0.0694277174836166,0.0515246050545974,0.0586726837070202,0.0030313890530711,0.00581214160453758,0.0925587774291272,0.0799999114309353,0.00891578533137238,0.00972978201500774
"1160",-0.0441778573307083,-0.0696571940689592,-0.0459999048587276,-0.053000857294477,0.0297531395682089,0.0132218610295127,-0.0235120859180827,-0.0527913921130917,0.0354071583215281,0.00428252295001075
"1161",0.0448836314686254,0.0488170940584871,0.0377358691599714,0.0552009447594457,-0.05044954636966,-0.0146924192854164,0.0466278156856716,0.0469799447211732,-0.0219383775697288,0.0216773984576242
"1162",0.00673359735104118,0.025128598087421,-0.00909093575931941,-0.00048476170167211,0.0198033908504511,0.00696503800438908,-0.00146103148019949,0.007803713053393,-0.00456807613469989,-0.00139135691917081
"1163",0.0211644403675313,0.0239551214696712,0.0122325310604747,0.0232615869712363,-0.0101351787103463,-0.00370149353352323,0.035655438751778,0.0210176197922187,0.0107666175750627,0.0121908874330814
"1164",-0.00853881031810388,-0.0174100231755671,-0.00805647944012156,-0.0085246032498919,0.0165547094893399,0.00459567195942445,-0.00370728922556196,-0.00839618592784985,0.0123399008322485,0
"1165",0.00066892800793994,0.0066444294641328,0.00101531657954856,0.00716477796238846,0.0175091439151076,0.00700818782259183,0.00124022744220431,0.00655549446827286,0.00287488503765965,0.00860291493408494
"1166",-0.0431184286802669,-0.0539054904104053,-0.0344828926883376,-0.0471895288502195,0.0205382207282081,0.00522048512939799,-0.0430091959230853,-0.033107272244328,0.0189198660580194,-0.0245650104809031
"1167",-0.0163307258575126,-0.020057913364081,-0.00945371819301777,-0.0124444152088452,0.0080682417480562,0.00105749703619429,-0.0199739522977326,-0.0117879736989015,0.0125478054661952,0.0178383776501641
"1168",0.000799285415011841,0.0115690345991322,0.00212092091829419,-0.00100790757279789,-0.00251791597123241,-0.00182479559618953,0.00188716277896139,0.00369225056505118,0.025784935133953,0.00171818966189541
"1169",0.0329103721196653,0.0340177354991213,0.0190474589476644,0.0350656793041195,-0.0137939194426033,-0.00404234248559843,0.024675223427741,0.0271650885139418,-0.0374884779779724,0.0102917024523768
"1170",0.0140843701659052,0.00425424121746221,-0.0114225752084994,-0.00974914076928501,-0.0284306056185787,-0.0107255347765844,0.0112133547899096,-0.00110243106996089,-0.033883064489031,-0.0101868622966957
"1171",-0.015244191364823,-0.0276761402479556,-0.013655428346066,-0.0194435956443705,0.0108211739421558,0.00615390349775558,-0.0210869812328929,-0.0170984243279065,0.00413636484018753,0.0044597718600301
"1172",0.014534493682109,0.0116181805061728,0.021299341382919,0.0170683709112076,0.00986668456958495,0.00320345867765393,0.0148557935338212,0.0134677805397374,0.029647249769974,0.0112705134484055
"1173",0.0287357821942318,0.0267008723470199,0.0135556612181262,0.0323295301966693,-0.0138261134049671,-0.00657991185953666,0.0318393585042211,0.0271318277625823,-0.0201724346640422,0.00337722592734591
"1174",0.00263683735956866,-0.00782975197456015,-0.00411528511079129,0.00143437269706537,0.0160762119426903,0.00691541593436229,0.00390127276223362,0,0.0299615103223965,0.0134635385750419
"1175",0.00443778388545391,0.0194474247344436,0.0175621003175708,0.020530011097587,-0.0154540084327026,-0.00357944353831396,0.0107756193693693,0.015094320432639,-0.00770522028904908,0.00166055506291896
"1176",-0.0104725794972136,-0.010229576791546,-0.00913720056438561,-0.0053799996714442,0.0211986017000307,0.00796934353742995,-0.0167776281572817,-0.00929395232841645,0.000843990542178652,-0.00696293982860552
"1177",-0.0255502261482701,-0.0270947114029111,-0.0163931426234475,-0.0225776214802097,0.0324857806204053,0.00917053711549709,-0.0241734165859432,-0.0144730503564647,0.0301906457016543,-0.0053421641792456
"1178",-0.00729745162386519,-0.0422051026874712,-0.0218751715854105,-0.0103467906108388,0.010398888020182,0.00133917686815432,-0.00218567402329806,-0.0190375963880636,-0.00185555004760019,-0.00335688875632811
"1179",0.0282076553219297,0.0305755228513236,0.019169045380705,0.0296621656313032,-0.0190886604698763,-0.0053496456605755,0.0335886922004827,0.0202389439546462,-0.0318206243352855,0.00909395082323083
"1180",-0.0103912463609109,-0.0206516970327912,-0.0125388511379498,-0.0221961759374147,0.00896798317774117,0.00489836236785224,-0.00724104558388261,-0.018750002190943,0.0267110681419576,-0.00667547638088173
"1181",-0.0262099314407035,-0.0380158600728187,-0.0232803539460531,-0.0338081006680611,0.0106651310177639,0.00487413327530795,-0.0281089076891954,-0.0288011258354386,-0.00610528030477187,-0.0157930705888282
"1182",0.00646992525754908,-0.0101882741621309,0.00975077711455841,-0.00199943287636295,0.00105524419247538,-0.00304363702688892,0.00311180864572624,-0.00228067635220341,-0.0223021531096097,-0.0023899317720053
"1183",0.00917124213445808,0.00842151449492312,0.0171673132331831,0.0015027471958573,-0.014231190138307,-0.00295734360436251,0.000912337745673897,-0.00343024019976801,0.0105846777674159,-0.00308004014999508
"1184",0.0138438729271693,0.0238168696135812,0.00421934672025981,-0.00275096878863546,0.00846614852293448,0.000574838443595738,0.0056518292630594,-0.00372792880615092,-0.0074492329570105,-0.00480608216168577
"1185",0.01725737034063,0.0259820564362487,0.0115545580164431,0.0145437403726736,-0.0152880438048104,-0.00745976496474621,0.0193980447052671,0.0146803296699931,-0.0158569656847878,0.00413940847517402
"1186",0.00591846506661087,-0.00294462695921294,0.0103840934817514,0.00172984183647729,0.00726863883093598,0.00192724485783313,0.00818047915953413,0.0000858646125032614,0.00934635926650329,-0.00446586426941942
"1187",-0.00995681999006426,-0.031896309964725,-0.0143881898717412,-0.0296071917963435,0.0190665967608563,0.00817322974875445,-0.0197563896029523,-0.0234685300508576,-0.0154519173746062,-0.0169082305750911
"1188",-0.00116390226092145,0.00671162717036999,-0.00104269192158901,-0.0073734037490002,0.0041969463041347,0.00133569658998356,-0.0028794103545684,-0.00175869320279542,0.014251924461969,-0.00175497785306811
"1189",-0.0294583255916331,-0.0300001542222585,-0.0125262422928328,-0.0371419058080482,0.0330831812611272,0.00428667148072637,-0.0478253545336818,-0.025836717303435,-0.0124587723999247,-0.014767839573728
"1190",-0.0323243635885589,-0.0390501218537099,-0.0158560789070251,-0.0702312055244805,0.0375864651574009,0.00929505759134641,-0.0252082843087668,-0.0334539188494462,-0.0261535405531089,-0.0353319713791268
"1191",0.00602518210825376,0.0117033969500844,0.00322205941223008,0.0266096540171161,-0.0185993611033727,-0.00826955872744051,0.00803845910487544,0.00904280358706067,-0.054717538218559,-0.0177581084843996
"1192",0.0237800116772009,0.0285989004879224,0.00535344260199055,0.0150498096290106,-0.0160558912708937,-0.00416999488340886,0.0126729831014127,0.0117429365371935,-0.0138923714538353,0.00338990068006195
"1193",0.0111839089302335,0.0296782560967828,0.0159744364479735,0.0318508026066362,-0.0153082929836922,-0.00666077454031477,0.0105891290973037,0.018631663557289,0.0193552669202277,0.0168919313092548
"1194",-0.0204187728105326,-0.0182037220217237,0,-0.0300692027397691,-0.000341630963695994,0.000191764785651305,-0.0249570430261914,-0.0194904705598089,-0.0274544223540304,-0.0269472233298083
"1195",0.00790376625213884,0.0222495950741481,0.0178195798477347,0.0137174107368587,0.00692140018366105,0,0.0148494674683752,0.0149849635709332,0.00947379330768272,0.0117601987558278
"1196",-0.0249892730140706,-0.036577928051762,-0.0257465294477122,-0.0500678463680964,0.0251189473143523,0.00632182310001772,-0.0263767690860899,-0.0343478689436033,0.00228282185699724,-0.0344957184688444
"1197",-0.0284580054314562,-0.0313774893698094,-0.0158560789070251,-0.0210824883984602,0.0275199322806816,0.00925993149453586,-0.0470633627067012,-0.019032983989714,0.0183475201612997,-0.00504847487959281
"1198",0.0219230926486198,0.0223518385134995,0.0128892358665718,0.0154250954897528,-0.012681030916549,-0.00510304649612092,0.0377670484991444,0.0104964800603173,-0.0206262913495028,-0.001951653922452
"1199",0.0185153268641842,0.018694603747021,-0.00424181103924126,0.0232157268488773,-0.00719903300487412,-0.00417883513445749,-0.00759829953959779,0.00629522053419351,0.0115453438946038,0.0140790482234632
"1200",0.0180912532159154,0.0339035146065214,0.00425988064799987,0.0330532860518267,-0.018457414210153,-0.00696250995852965,0.0276043760189351,0.0272131655811345,0.00645928731208456,0.0208252518572627
"1201",-0.00669580454074781,-0.00842373571149124,-0.00530222530236757,-0.0119308446240792,-0.00738742151037153,-0.00518625511572413,-0.028235268747677,-0.0024360138180457,-0.00816257685330624,-0.00453344997004712
"1202",0.0334456109675239,0.0445993610862805,0.0255867485223,0.0447310806580383,-0.0141236274352218,-0.0105227656681623,0.0482242819449217,0.0335777035824913,0.0256942529203403,0.0223909381486429
"1203",0.00100341055185149,0.000290655908433468,-0.00831642518880771,0.00052550686147379,-0.00334589459396806,0.00331690245635308,-0.0184792825702049,-0.00797436851253019,-0.00716603155102513,0.00742391804903431
"1204",0.00877195071374426,0.0223577428801638,0.00628948910641092,0.0280914492962883,-0.0145463621062274,-0.0034036148083546,0.0162778242822401,0.0214352227888961,0.00715600837177011,0.00184234981324116
"1205",-0.00198744601398859,-0.00198810702893648,0,-0.00893792736060706,0.00995737576605271,0.00400055309500247,-0.00694728026255542,0.00466319363363299,-0.00588014228470357,0.00220658761071491
"1206",0.0170938500712083,0.0133750548698148,0.00208357440374507,0.0200981036376631,-0.0145296077879585,-0.00495646407381678,0.0231248462885978,0.0165359942384478,0.00677751681865324,0.0227523610500662
"1207",-0.0190910626148514,-0.0292051614887662,-0.00415827297254789,-0.033847007027768,0.0172885096025805,0.00654407888235942,-0.0229821936390926,-0.023116253255955,-0.00477355586683803,-0.0143524120639776
"1208",0.0195458153004309,0.0161989258215751,0.00939471961353777,0.0266668701751487,-0.0062109761554997,-0.00106693719143724,0.0330482817946121,0.00964056112082967,-0.00479645199841494,0.00546057776377684
"1209",-0.011828885889984,-0.0170793784321085,-0.0155122139621519,-0.0190988112247849,-0.000346701684626582,0.00155381233527807,-0.0124201938064149,-0.0144676930302475,-0.0121725225450452,-0.019551117232251
"1210",0.00437560151314775,-0.000868722365076957,-0.00315122922893984,-0.0192107404994942,-0.00712086990863359,-0.00203699342862029,0.00609781295496159,-0.00411050308616201,-0.013135616849178,-0.00147700870732781
"1211",0.0189872178207136,0.031594107422817,0.0105374967033312,0.0285865610740714,-0.0105827491148728,-0.00184610544048447,0.0295455456012881,0.0250593912642778,0.0110920958080218,0.00517744365051964
"1212",0.0122607962747614,0.0126439060770756,0.0104274037522314,0.0391146794649668,0.0016795577398816,-0.000486870738336531,0.0264900422994665,0.013229796660267,0.00940320939309913,0.0158204292876116
"1213",-0.019444026726174,-0.0174803820301189,-0.0144477910397794,-0.0198118182308182,0.0254144936227942,0.00857244041957572,-0.0154126770081029,-0.0218565858438923,0.0283815171188295,0.0032597558763543
"1214",0.0101589079909679,0.0180739569148176,0.00209390562313794,0.0184440500826031,-0.017469589640546,-0.00734075369192211,0.00928349944824114,0.0078352934050494,0.0109305999379332,-0.00577620555844283
"1215",0.0348351783455707,0.0590846111786982,0.0386629724874812,0.0607784680155465,-0.0338963123776266,-0.0120654001997673,0.0427410782182294,0.0457814971614527,0.0128435428737232,0.0265069102104287
"1216",-0.000233413802483873,-0.0125719271849242,0.00402385081605661,-0.00841894423264211,0.0105164979374366,0.00600816591356335,0.00311319177500535,-0.000825774369188625,0.000412810373114469,-0.0042447971617956
"1217",-0.0241056133773228,-0.0498676487960267,-0.0581160768172869,-0.0375000716546834,0.0396553487553659,0.013411956057608,-0.0131034945796399,-0.0338932740612079,-0.0134418056078823,-0.0152752847674487
"1218",-0.0278884349897368,-0.0424342470749794,-0.0127657986300936,-0.0242585524657136,0.0334744877558919,0.0119943660581403,-0.0337175675338868,-0.0199660208315005,0.000239088089855066,-0.0119047844473724
"1219",0.0163113438469309,0.0134108866221989,0.00323269441168872,0.0306377410726035,-0.0124736142224054,-0.00239117413242707,0.0202497972090929,0.00407438010070815,0.0100369993417075,0.00620655986768326
"1220",0.0182271466537181,0.0322209202246699,0.0075186689316642,0.010233916214238,-0.0137341285037325,-0.00469847827701997,0.0113409257368,0.0133331505036163,0.0157340768453103,0.0123368135976034
"1221",-0.00609879764092025,-0.0167223702217287,-0.00213231934793556,-0.00651223668070111,0.00120384880852087,0.00298656654530061,-0.00753456453520573,-0.00514898976830802,-0.00506635799518773,0.00322572541378996
"1222",0.00621622820797829,0.00113401910462474,0.00854710003886527,0.00849710709619633,0.00635270825702583,0.00115282714933573,0.00247172598099055,0.00373820918963474,0.0241731920103063,0.0146481467086375
"1223",0.0128305934259485,0.0181199747405378,-0.00423722543291438,0.0117960438598372,-0.0127967814820532,-0.00450937322524969,0.011975879106376,0.0117442541484596,-0.00828664437733784,0.00492958259453546
"1224",-0.03690960244074,-0.06312577326309,-0.0180850384454477,-0.0585300132447313,0.0207406020242988,0.00886655695074845,-0.0449006297059032,-0.0450164839804162,-0.0084134847485362,-0.0220743406300569
"1225",0.00941870274852641,0.0175127448804173,-0.00108345464014614,0.00657098615474427,-0.0149007524700291,-0.00487238713105365,0.000911200812269142,0.00326082372769387,-0.00540482339842074,-0.0010748689279797
"1226",0.0188222540549496,0.0306298851318718,0.0108459828851883,0.0241024508480532,-0.00610166393526745,-0.00460749533401772,0.0258508107611157,0.0260047779289776,0.0164777843664707,0.00968441420898558
"1227",-0.00947409626925844,-0.0209451081649991,-0.00429171924537941,-0.0137290209315415,0.0160832493445484,0.006269211779804,-0.0200531955426234,-0.0207374956177951,-0.00436887772716632,-0.0106571575633633
"1228",0.00494165796390811,-0.00578214179349423,0,0.00621450724461159,-0.00136161799350121,-0.00134258377391505,0.00869268281480506,0,0.000923810639557932,0.00718126704142441
"1229",-0.0158631309757555,-0.0180284590440442,-0.0183192067056729,-0.026926985845745,0.00911808465608299,0.00364742754445602,-0.00951528052522499,-0.026764762041125,-0.0106714697123242,-0.00249550960909894
"1230",-0.0158763972863994,-0.0106604779922673,0.00109775831917358,-0.0253870431939014,0.00802232516908474,0.00200791333841766,-0.0179443859559684,-0.0163188553970252,-0.0257127230398438,-0.0232309291562415
"1231",-0.00106490466687126,0.00329247516761644,0.00438602720397907,0.00390701616493927,-0.000251102923569668,-0.00372193704187296,0.00719796401134509,0.0061442682653603,0.00311184309592405,-0.00146353550983858
"1232",-0.019019409536202,-0.0256563086998787,-0.0196510280070411,-0.0321742357403266,0.00594913977621703,0.00277798524832273,-0.0263882852199321,-0.0262592990551541,-0.0245793767026421,-0.00732866692535983
"1233",-0.00392791491228417,-0.00979796109185027,0.00779542362925922,0.00348522736363055,0.0111621370625445,0.00305623523712328,-0.00282306178664216,0.00689838771668305,0.0110703241590215,0.00664450312592546
"1234",-0.0220653381317847,-0.0303029248750388,-0.0232042840811086,-0.0323268607345555,0.00980272388967474,0.00342829995046245,-0.0294451648304832,-0.027717129183745,-0.00290361143189899,-0.0150348950280789
"1235",-0.00188782616641003,-0.00510212553172085,0,-0.00331331190169459,-0.014521022624793,-0.00635822748334736,0.00350097653865578,-0.000640617384381814,-0.00867565359854827,-0.00819058292561925
"1236",0.0289672981564315,0.0503205428053579,0.0282803000093368,0.0479227823289705,-0.00049697860555098,0.0000954682040517074,0.0244180749376826,0.0326922250429482,0.0197675099057839,0.012387333873749
"1237",0.00283985833924083,0.0064081749834326,0.00440069465415593,-0.0044939181234025,-0.00819924508642966,-0.00191028956986716,-0.0028375877112915,0.00682803358356998,0.0015003300275962,0.0129774726077585
"1238",0.0411494416972424,0.0527595038504769,0.032858532832799,0.0624002711272944,-0.0156157605366971,-0.00583613137017103,0.0461014308924579,0.0554871184468333,0.0194750713244525,0.0117129078004778
"1239",-0.000159679060676821,-0.00576064294195378,-0.0137857549888084,-0.00299914931454448,-0.00501814514096199,-0.000289851446918621,-0.0101559642312153,-0.0175232907081708,-0.00293892896787962,-0.00361785859813823
"1240",-0.000880319187381962,-0.00144831555526681,0.00322577411568137,-0.0030083243616158,0.0140182282139845,0.00443693364212683,0.00164890937223383,-0.00356714763590893,0.00112009664799562,0.00871458986637008
"1241",0.0108920675543476,0.0104440670863994,0.00750270832044775,0.0163439724904557,-0.00202331002567402,-0.000575664503775442,0.00932875449120285,0.0137231530605906,-0.0147214691847233,-0.00539956831462385
"1242",0.000317122642589096,-0.000574297531647505,-0.0117023090563975,-0.0136071277497335,-0.00954372430379424,-0.00259446262566598,-0.000724911042369158,-0.00706309820213413,0.00513976789398529,0.00542888193349578
"1243",0.00372243777121795,0.00660722071049502,0.0139937580853877,0.00401318295601927,0.00358150638706056,0.0045278390287613,0.00943055275214966,0.00533474479085294,0.00725413872505043,-0.00863930189363515
"1244",-0.0219363194458232,-0.0342466415784847,-0.024416280998294,-0.0359729937784271,0.0124902339096122,0.00508345441422442,-0.0238952603400027,-0.0341977773861811,-0.0201888909157812,-0.0127087255023969
"1245",0.0169420020981348,0.0257094201930046,0.0228510462700369,0.0202122651818049,-0.0205604399497192,-0.0068705339241244,0.0198788435369566,0.0149571238126442,0.00253041336378867,0.00367777219365739
"1246",-0.0145971637620048,-0.0342842223026918,-0.0170215179761157,-0.0375919591458623,0.0111389726522528,0.00345894723511053,-0.0178669652333903,-0.0315787292976352,-0.0265023386959977,-0.0128252236904338
"1247",-0.0093395276016518,-0.0167065080028356,-0.00432890962891586,-0.0092372200249129,0.00932092211834501,0.00459596434773357,-0.00882018528444151,-0.0102485329546853,-0.021853249526105,0.00408313009436156
"1248",-0.0106457909989298,-0.010922542825796,-0.0108692790530927,-0.014384739706484,0.0188900264496377,0.00419293325269265,0.00574704841725415,-0.0128651104381142,-0.0350899217751327,-0.0354898435017028
"1249",0.00361439786341666,0.00429487746227153,-0.00219805645903681,0.00648649894107201,-0.00370806093544507,-0.000853881439196735,0.0136403538633272,0.00985397403147381,-0.00366274448075565,-0.00498276289883115
"1250",0.00148232054095643,-0.00763592350234132,-0.00330386806456295,0.00751877307267113,0.011661667869677,0.00484431535327445,0.00836557598161791,-0.00331912797469647,0.0190375760646284,0.00808941651852191
"1251",-0.0106913316609266,-0.00447576447369147,-0.0143647325457791,-0.0258527480031721,0.0126720007226457,0.00340395237374769,-0.00973863235299288,-0.0150495383328703,-0.00231914584343618,-0.00458549768908145
"1252",0.030259985398351,0.0384012878374869,0.0256409379843743,0.0419025155577646,-0.024945653883527,-0.00904514025732117,0.0302310292943193,0.0367361479680481,0.0136243369801878,0.0230327116103957
"1253",0.001936839981588,-0.005411591615607,-0.00995578504519667,0.00318127109789068,-0.0139097159862281,-0.00323261463296498,0.00141449583224396,-0.0119161811199424,0.00114669387556865,0.00712943567986613
"1254",0.00885854132415598,0.0120918880092367,0.00670405051147616,0.0132136236106333,0.00419815374933985,0.0012399849826219,0.0136807903411116,0.0111077160918112,-0.00712656510240339,0.00111779615846253
"1255",0.00894082064133284,0.00567500568851109,0.00776912064933599,0.00391217250969289,-0.011120445096552,-0.00409606822218778,0.00492685457831277,0.00784668123746779,0.00173035767823948,0.00483808137586306
"1256",0.000790996306225367,-0.00267305818011099,-0.0121145939708436,-0.00961288525545034,0.0047504660046287,0.000565394730420277,0.00227641403689893,-0.00653997823345376,-0.00895652241003819,0.00444445986150788
"1257",-0.013123180477069,-0.0157831728182188,-0.0122630931564852,-0.0167890849621181,0.0184883715031274,0.00632149266509541,-0.0108315482539918,-0.0163008389480789,-0.0250468329985969,-0.0117995140293872
"1258",0.0103339137342271,0.0160362761358313,0.020315996307378,0.0114729776715849,0.00182363050554768,0.00123675011397695,0.00830114175331942,0.0114723031879587,-0.00456864864310824,0.0029851108523391
"1259",-0.00491597597760596,0.00476477582265478,0.00774346596550002,0.000791283853265101,0.00322666863118815,0.00351744554575517,-0.00490487762803771,0.00283547106513393,0.0109751832107272,-0.00148807495388825
"1260",0.0159361907838804,0.0314166139318277,0.0197584127723933,0.0305745836608611,-0.0150098444211564,-0.00634646072368994,0.00616103652014943,0.0248192462377828,0.0258569173676915,0.0298061975373973
"1261",0.00156865122737937,-0.0103448202686788,-0.00107608315000385,-0.00562665895381165,-0.0118899426861534,-0.00314594804820822,-0.0111966373705679,-0.00367836369667029,0.00506675865914263,0.0075978046715317
"1262",0.00266245750357896,-0.0185830296909629,-0.0118536549751319,-0.00437261386086973,-0.00177979326251243,0.000191430617863642,0.00725415217302183,-0.0101540706761304,0.006827847311627,-0.0136445958527361
"1263",-0.00257726906704736,-0.0121303028389966,-0.0109051841410253,-0.0126580715868017,0.0078949949111502,0.00392003641626726,-0.00175664451513313,-0.00590603738773765,-0.00367601726249223,0.00436834231689986
"1264",0.00242749356572713,0.00509147745776284,0.0033077868676239,0.0104655648304606,-0.00176891614885633,0.000190040197847852,-0.00281525473992983,0.00250120242059415,-0.00445290720966107,0.00108748494039279
"1265",0.00867055503785785,0.0146008395453785,0.0120879662863933,0.0217504510499731,-0.00168736622381271,-0.0019994107200908,0.0111167498191005,0.0155960569717657,0.0136741150159743,0.0072410675824528
"1266",0.000541954943797496,-0.00616752877450166,-0.00434327751971086,0.000760539435749497,0.0130159369271539,0.00582029189755162,0.0089007797031464,-0.00061434354197365,0.00649268158404359,-0.00287566377870796
"1267",0.00239922091784806,0.0100472357295183,-0.00436191092656435,0.00405174918729267,-0.0014183301943318,-0.00208731501794668,-0.00657340563917053,0.0129070620517204,0.00444671515559247,-0.014059040274147
"1268",-0.00517333786727392,-0.0184317241424796,0.00219047884267942,-0.00907947177799062,0.00994184934772568,0.00446780204293296,0.00452716898464045,-0.00697811262311832,-0.00698347652501952,-0.00219379185917579
"1269",0.00388074877830169,0.0157972856225548,0,0.0190887882416446,0.00463320074661522,0.000946051264288261,0.00520031649057384,0.00824950250529266,0.00778604193727372,0.00696219963645928
"1270",0.011056239098624,0.0184858444136229,0.0120216618986624,0.0252246452224361,-0.0121050501293039,-0.00311963828370321,0.00638039839420079,0.0139391620854561,0.00685361993769473,0.000363970964420313
"1271",0.00527661284277303,0.0164218251160504,0.00755968195654821,0.00876982033858464,-0.0137535067274204,-0.00597494213516625,0.00633987564311478,0.0197253009046809,-0.00235151600180017,0.00436516390143638
"1272",0.00372731818365257,0.00255107361904616,0.0128616624569855,-0.000724725430670037,-0.0113254652801372,-0.00343447467687674,0.00476765305715787,0.00820600109046232,0.00527233590576648,-0.00724372798843753
"1273",-0.00257691913543867,0.00763356345975863,0.00423269924987224,0.00966659326546515,-0.00632525388032379,-0.00220205029913556,0.00305037500431982,0.00668637264833682,0.00672547018523906,0.0116745244053
"1274",-0.00113949412254688,-0.00280561588483375,-0.00948357642845565,0.00143615161172117,0.00180590514538848,0.00115110565962628,0.00557556227169953,-0.00779674940776742,-0.00704835113879987,0.00180315100471051
"1275",0.00836750798530828,0.00675258322744576,0.0127658852176988,0.0112334414603301,-0.00240391918773708,0.0047921791217227,0.0127684033098039,0.0130964034424617,0.0272205612993197,0.00827933561250238
"1276",-0.00512969817777542,0.00251575037087926,-0.00210095419818568,-0.00401796139283583,0.0132563300051443,0.00534133792624369,0.00580637778278459,-0.00229785914877367,0.00510759530233873,0.00285608377297009
"1277",-0.00045501844225293,0.000557387850526947,0.00526329271398884,0.00522054773736391,0.00314329875622632,0.0030358506603354,0.00247422281954335,0.0051827602543002,0.0101631910046465,0.00356001051713029
"1278",-0.00341408757109785,-0.0153247529512519,-0.00628276241059234,-0.014400289569131,0.0117717804467725,0.00340551498658703,-0.00872006188905528,-0.00773398889106869,-0.00556312951670035,-0.0102873049938557
"1279",-0.000380228161096396,0.00679142362024954,0.00632248508220834,0.00862278121893056,0.011550900921961,0.00377075682032246,0.00514511682452312,0.00346390750536041,0.00761768141175789,-0.00250900001479271
"1280",0.00875722023667347,0.0207978909964619,0.00628285255755334,0.0220850090909781,-0.0114553582971542,-0.00347211578618545,0.00743069799573348,0.0161103256402333,0.00147658143614171,0.00323395006293814
"1281",0.00158502499006863,0.00220299855077521,0.00312176759974792,0.00278824384626941,-0.000418941633091863,0.00141657783235716,0.00213080507742469,-0.00141544136925964,0.00878747946198954,0.00250709217230694
"1282",0.0140186788346832,0.0189558655702915,0.00311205249510005,0.0166818537837308,-0.0214895653182604,-0.00791951470009711,0.0143930132916048,0.0144597897988905,-0.019935714353656,0.0117899484229973
"1283",-0.000668727080547327,-0.00620100524875367,-0.00310239767068821,-0.00843214125670011,0.00995122455231057,0.00275615031174148,-0.00483716052394056,-0.00614842794870052,-0.00274401099226917,0.00494350813762146
"1284",0.0025285232340535,0.00678225559927625,0.0103733793204168,0.00206860099034167,-0.0124008514123881,-0.00644445248842129,-0.000810145801952045,0.00337415739152735,0.0150735979514007,-0.000702731107745658
"1285",0.00296774008774903,0.00323373205846034,0.00410679209182718,0.00711006241771583,0.000774290597976846,0.000476768550004447,0.000648925775380338,0.00532534494775883,-0.00707128474492547,0.00457096435919468
"1286",0.00125757577793584,0.00268614281737189,-0.00306750383408627,-0.000455724985551575,-0.00747698670672947,-0.00228793713536979,-0.0072922217898157,0.00139386979413114,-0.00284864094955495,0.00525029928143272
"1287",-0.00738758021092367,-0.0192877296574149,-0.0123078577641582,-0.0221003216364338,0.0129883236570048,0.00563774759591373,-0.008325408726924,-0.0153120596600197,-0.00523750136323065,-0.00940102202020787
"1288",0.00744256274014132,0.0101065036021653,0.0103840345033694,0.0163092100374984,0.00128188498475801,-0.000664816016026415,0.0113581495589175,0.00706849571961343,0.00221368913613551,0.00246042320711748
"1289",-0.00125599626745276,-0.00892343882738178,-0.00308291416996476,-0.00825312150052471,0.00529261088951394,0.00209143373066589,-0.00992844585837838,-0.005614964612633,-0.00232821928028837,-0.000350626340403282
"1290",-0.00466001445473962,-0.00300155576522187,0.0164947911940883,0.00277386886331499,-0.00178293693003884,0.000759306725986564,-0.00493162857441631,0.00847018371171182,0.00592392310686707,0.00350749322354549
"1291",0.0110727457361304,0.0139573139017426,0.0101418095439967,0.0108345411096187,-0.00799663753475133,-0.00455079894272548,0.00826029262032901,0.00895828708079205,-0.000654339416725214,0.00454391175146429
"1292",0.0026465029883167,0.00431831028813612,0.00100412824605756,0.00182429081122337,-0.000257586574435087,-0.0010481542754478,0.00163863302379297,0.00721433594939103,-0.00386901190476185,-0.00173971176077381
"1293",0.000439837808570598,0.00134377621380333,-0.00100312098394351,-0.00409723495504521,-0.011065082592302,-0.00362322662922421,-0.0124328241473344,-0.00688726862301692,0.0219300739074966,0.01568487205973
"1294",-0.00322426354565042,-0.00509914235990983,0.00301238473817267,0.00182868168260297,0.0125765246192218,0.00392420503334612,-0.00811620380774913,-0.00693459480263059,0.0112267451473103,0.00926559358588586
"1295",0.00441070065531601,0.00971110426794874,0.00600569839296039,-0.00182534370999599,0,0.00142944018011693,0.0116899774406181,0.00810024240405793,0.000462599740226777,0.00306014184494452
"1296",0.00219560467061974,0.00854942558352167,0.00199018638434278,0.0100570579544599,0.00651060124296077,0.000760929586009373,0.00280593519780159,0.0119146722982493,-0.00456599226526433,0.00610175144674652
"1297",0.00167996410588223,-0.00741741924576689,-0.00595790230452542,-0.00995692062666953,0.00885103891318573,0.00332907841129204,-0.00115217238047272,-0.0049288190870076,-0.00307727464616558,-0.00808621224280259
"1298",0.00291639853022385,0.00854071441073367,0.0159836428977225,0.0139431033119706,-0.00329004710049374,0.000474254892986137,-0.0075808646380654,0.00963154842209701,0.0104252069381223,-0.000339669258072273
"1299",-0.00392567263401156,-0.0108496082828715,-0.0176989729599565,-0.000676339189776165,-0.00609392579882218,-0.00397980948369325,-0.00132843317272247,-0.00572393747541766,-0.0530290606654832,-0.0037377712839286
"1300",0.00518186309015967,0.0136435612391028,0.00600569839296039,0.00947428379056059,-0.00941437666835643,-0.00323982945694146,0.0053212396104434,0.00986862018593659,0.0141214200429116,0.0156890517662007
"1301",-0.00304958231587449,-0.011348649167926,-0.00995018951728954,-0.00245823506448717,0.00939178071788893,0.00401555178725754,-0.000330921880576818,-0.00488583439199708,-0.00162058098781237,-0.0100739096678047
"1302",-0.00407819655551822,-0.00400404336752747,-0.00602992991005014,-0.0172488847998162,-0.0079384041132281,-0.0019994884662613,0.00810723801177926,-0.00436457373686505,-0.00414814245877471,-0.00474902210510297
"1303",-0.0146252990283687,-0.0399358949962484,-0.00808912563585917,-0.0335082179596229,0.0121322763429919,0.00419748020015676,-0.0134580358806528,-0.0263014199585709,-0.0178086151937923,-0.0163598703524483
"1304",0.00697609446651315,0.014237935555407,0.00611621752301605,0.0120282991412197,-0.00612048805381282,-0.00190006586241509,0.00432507063797827,0.0123803390090007,0.00571609107036442,0.00450444281824036
"1305",0.00994887365288766,0.025323224636888,0.0172240006280144,0.0209742963331732,-0.0100084569970972,-0.00295079867235593,-0.00231873469241994,0.0216787079107188,0.0100836885019957,0.00827878144789507
"1306",0.00386724935823768,-0.00697958303362367,0.00398396478825114,-0.000456654671093792,0.00198722147627217,-0.000763495690851768,0.00464889281606906,-0.00516850103221667,0.00665540904317163,0.00273687664164446
"1307",0.000072846022603601,0.00162191840931158,-0.00992080228916059,-0.0109615697488147,-0.000171868491535609,-0.000286691041748721,0.00694095621642732,0.000546634278952185,-0.00787353023579973,-0.00136470329624794
"1308",0.018025883846517,0.0178135413546809,0.00901820986564505,0.0272458565629337,-0.0175945344553682,-0.00716744468676189,0.0178891753297259,0.0177645240002331,-0.0167807831982463,0.00444138199630006
"1309",-0.0010710114438508,-0.00689444412378282,-0.010923699558423,-0.0157341098078142,-0.0251952102219297,-0.0114544132972044,-0.00241845714995736,-0.00939835350402507,-0.0168206774463214,-0.00680273323384251
"1310",0.00578958229353277,0.00961284353694047,0.00803239210368134,0.00799260752801434,0.00153145988395265,-0.000291847114404553,-0.000646424072635932,0.00921653157667057,0.00946289987942417,0.000684922163946666
"1311",0.00138460144664587,0.00872779075040397,0.00597610438585128,-0.00113251254654856,0.00197783398755558,-0.000292630524992177,0.00598407064902706,0.00637943575600186,0.00136578716953339,0.0123204071609913
"1312",0.00392002041516859,0.00471945079320424,0.00296997461641979,-0.00385585777113007,-0.0119354976831867,-0.00613789174003154,0.00594838528013342,-0.00134293750382586,0.00179784869563826,-0.00169030813224702
"1313",-0.00291074322303342,-0.011743256217028,-0.00987180864018089,-0.0173040740124243,0.00399622626567253,0.000490170502587706,-0.00239719862078769,-0.00995192692913449,-0.00903515710217606,-0.0121910687751201
"1314",-0.00163736226408573,-0.00580941171978833,-0.00498485893695244,0.00185334309935636,0.0113080995320731,0.00509478515548234,-0.00224293816648569,-0.00353153744722812,0.000499606554061893,-0.00239976354492633
"1315",-0.00720399688714723,-0.0114209230619514,0.00100234600550508,-0.01526361380588,0.00322040918973898,0.00126751778464085,-0.0118818246576299,-0.0109047238658622,-0.00399475670705129,-0.00790370781297056
"1316",0.00323273906423216,0.00698531227714683,0,0.00751523526282449,0.00945173782537556,0.00369990228620432,0.00406262211248332,0.00303173007033819,0.0122829599173986,0.00969855199605174
"1317",0.014035284089126,0.0170757637114787,0.00700704070699665,0.017482598631116,-0.00512323754501731,-0.00116410060070782,0.0103333255596418,0.0129157212538107,0.0177675665063304,0.0044597718600301
"1318",-0.00310707804224553,-0.0115422527980634,0.00795220200978974,-0.00526924068279511,0.00719162503255233,0.00553570252855695,-0.000484800370922023,-0.00189922284625499,-0.00705589441809829,-0.00409837491775156
"1319",-0.00495845177021881,-0.0111466595368095,0.00197240830162171,-0.0168124971789569,-0.00141040260407044,-0.00173852207974101,-0.00226316535143523,-0.00679516438070105,-0.0105979536082469,-0.00960224010502808
"1320",-0.00170900883510572,-0.00778308816498408,-0.000984474619182274,-0.00117095079646046,0.00750328002584233,0.00416014094757355,0.000972182248560438,-0.00191585530905181,-0.00142403570751148,-0.0138504051469359
"1321",0.00413640295706519,0.0102785618452084,0.00295588193051377,0.00726979610280742,-0.0169103925501157,-0.00491388234092072,0.00841705466175657,0.00959706301809837,0.00520830856403953,0.0112359826673936
"1322",0.00731475907447821,0.0152611205733526,0.000982004892828847,0.0137370982237972,0.00553970457228914,0.00239580785738402,0.00642062496259688,0.0103204591230508,0.00505802507580877,0.0128472255229006
"1323",-0.00408926569997914,-0.020833232257916,-0.0127572287531899,-0.005741927859927,-0.0173283278813867,-0.0073536818479768,-0.00462535593696556,-0.0129032445497825,-0.0187185648862335,-0.00445657267375199
"1324",-0.00991052008922444,-0.0258552909462586,-0.0228631441591989,-0.0180181527118458,0.0137455586218511,0.00506893784283413,-0.0100945479019438,-0.0152506879607111,-0.0167614736178715,-0.0154959387610798
"1325",-0.00050086469330346,-0.0091236665825748,0,0.00541057625492947,0.00722596073723736,0.00446108502316744,-0.00437045974123929,-0.00359497522133168,0.00699695280848123,0.0038475546290011
"1326",-0.0112307576224931,-0.00446417468456195,-0.0061036575207023,-0.0147402301776123,0.0233812969396525,0.0102348390743687,-0.00959194581923983,-0.00499600167714376,0.00669570471474579,-0.00452973397957102
"1327",-0.0167851698387155,-0.0252243067780112,-0.0122826637241058,-0.0194726600700478,0.0113372858534317,0.00468318029335912,-0.0193693231379809,-0.010878534039191,0.0108553118797552,-0.0133005924675427
"1328",0.00809442042243047,0.0169639670524362,0.0134717888420761,0.0108984299565351,-0.0119803168811141,-0.00390075244764199,0.0118844137353151,0.0118442665437899,-0.000186213525032453,0.0024831161464689
"1329",0.0130660521935069,0.0197907675636171,0.00511225209011901,0.0256346128385194,-0.00415711486060422,-0.00200481806158448,0.0142268518082145,0.013935490911869,0.0101197611545394,0.0130927143080344
"1330",-0.0118889377885906,-0.0263376743596981,-0.0111901701567613,-0.0151832257888399,0.0161770164276243,0.00602833251167589,-0.00521936086343611,-0.00769643620268168,-0.011370565667558,-0.0101291689588564
"1331",-0.000656041002875085,0.0105351333490462,0.0020577542859106,-0.00498096613480192,-0.00145514580771389,-0.000285550017496305,0.0116412941957245,0.00332378952008616,-0.00242461290302975,-0.00988007454080853
"1332",0.0148122108802209,0.0208510043798458,0.00615984931538738,0.0114420455948054,-0.000600174660627451,-0.00104629630363462,0.00858988679144268,0.0124241195463015,-0.00130878094751663,0.00463293958054045
"1333",-0.00337946193480676,-0.00800417849371682,-0.00204048812418534,-0.00471367384545263,0.00291565539063421,0.00200006261893448,-0.00530289365276071,0.00245416869749837,-0.00586584711388449,-0.00957784323772171
"1334",-0.00642095291357281,-0.00528707065103884,-0.00613512503741498,-0.00449897015875345,0.000941063583635104,0.0011411054899646,-0.000484655337972373,-0.00435246523375177,0.000753217007761098,0.000358161290763714
"1335",0.00167015839659257,0.0125877153833478,0.0020577542859106,0.00689821879107422,0.000170732573600896,0.0000944137944300927,0.0105059796691296,0.00928968796919172,0.000689958005580582,0.00393840047884164
"1336",-0.0084089376774148,-0.0223757282759129,-0.0112938034694821,-0.0191356156432166,0.00726051592396648,0.00199352903322647,-0.00927719185938425,-0.0143475875540182,-0.00294588203974666,-0.00178321596697351
"1337",0.00380139039193161,0.0073467397428375,0.00623056969882918,0.00216774641696693,-0.00703878146906234,-0.00255827765706629,0.0127544164080751,0.0120842704836495,0.00144587910906413,0
"1338",0.0136915744830985,0.0165497597221038,0.00516009044373411,0.00913244730683838,-0.00512404244887055,-0.001234972946763,0.0109994063322816,0.0108551418662413,0.00200873819192582,0.00571639657127987
"1339",0.0069688929106797,0.00662269080897482,0.00513336489782734,0.00619197784824443,0.00600894553905551,0.00332923413154163,0.00425744261997685,0.00375842490947997,0.00883350485006607,0.00213140957556313
"1340",0.00164095599586855,0.00520816907643074,-0.00306445883758633,0.00142017524466587,0.000853299445335853,0.00104233897810624,0.00486728789380253,0.00401186560463862,0.00217354531561553,0.00319035098056442
"1341",-0.0037037259924575,-0.00627199376591636,-0.00204896818440803,-0.00212715603150138,0.00025573880360219,0.000852493296819246,-0.00140645128104211,-0.00372955712406198,0.00309827726179579,0.00388694552119162
"1342",0.00621998846653282,0.00768371511326893,-0.0102668771097216,0.00663141013270185,-0.00518616904595692,-0.00181972881067927,0.00876241508851816,0.00267370866547023,-0.00345934014518967,0
"1343",-0.00298423339969123,-0.0106207840478448,-0.00518673431287187,-0.00188223945505128,0.00704307768764201,0.00189906397572415,-0.00155107505631669,-0.00239968303283378,-0.00452523536029847,-0.0130235865097412
"1344",-0.0076252973561528,-0.0090834123654745,-0.00834217452459174,-0.00754335547860563,-0.000256264076453183,-0.0000947532399543372,-0.00341758920985646,-0.00908858768791865,-0.0100877703490323,-0.0110556673761554
"1345",-0.0161581590926256,-0.0172223159323822,-0.00736058908128745,-0.0175770504403667,0.00784906332396473,0.00398040170345126,-0.0076386036238506,-0.0129486644129603,0.00314524751119549,-0.017670375073744
"1346",0.000729801818543541,0.0081967336179305,0.0042371830267296,0.00362666203972739,0.000168675936107254,-0.000283082174927785,0.00565518266280418,0.0081992483002169,-0.00244559476738193,-0.00220261312828607
"1347",-0.00401165543330417,-0.0134568578787305,-0.00843873120137417,-0.0158997494067412,0.0053316522615261,0.002265995401034,-0.000937169325562648,-0.0103011302766454,-0.0193613399627692,-0.00367920130409782
"1348",-0.00593169289798989,-0.0147768800132925,-0.00851067155444096,-0.0129744400542772,0.00067369956855079,0.000847831240932795,-0.00234522867862441,-0.0106819662951885,-0.00980768589743597,-0.00775473278825167
"1349",0.00206290926038677,0.00519195475525169,0.00429173924638127,0.00421626908223161,-0.00294464199819555,-0.00141210862724139,-0.000940339819027969,-0.00027674606298167,0.00194214409307869,0.000372080552337062
"1350",-0.00301450341287557,-0.00487798929870731,-0.0106838192502329,-0.0128425852668614,0.00826895325870391,0.00329939916607924,0.0042353177077652,-0.00498493350747164,-0.00781809115931786,-0.0074404513480204
"1351",-0.011060980377558,-0.0204729342515516,-0.0107989479869498,-0.0227671296387799,0.0139746084316423,0.00441539336781283,-0.0121834592043275,-0.0125244855554021,-0.0145219850810365,-0.0131184545155544
"1352",-0.00574161600242173,-0.0156019323590428,-0.0131006132965846,-0.00870467909331807,0.00404421339755867,0.000280513796449444,-0.00490209562841648,-0.00930053757599858,-0.0105068193946103,0.00189894864774565
"1353",-0.00382485478445427,-0.00687815891448995,-0.0110616271427159,-0.0142044191463745,0.00287686891806449,0.000748305286388362,-0.0122357092467047,-0.00825067382790357,-0.0018698944213339,-0.0011372096858524
"1354",-0.0148312279567023,-0.016561323935297,0.00894835491711898,-0.0136232930156444,0.0177035714699671,0.00373757953889386,-0.0276706088966919,-0.0117610648944485,0.0223470884756483,-0.00227693068930646
"1355",-0.00855873024948972,-0.00275568250675351,-0.0144123705403665,-0.00956184754100509,0.000241514176507529,-0.000652049753838591,-0.0102580034104613,-0.0072569485552938,0.0114528793562916,-0.000760813374248825
"1356",0.0171883327543956,0.0239485631387193,0.0101234110085373,0.0238671159152162,-0.00209327827047867,-0.00260760949965921,0.0205615412554765,0.0236839152499446,0.000646981546807091,0.0133231960579028
"1357",0.00174272982907842,-0.00329836775005621,-0.00111342269049475,-0.0104764652398107,-0.0111348704341897,-0.00214839401342071,0.00212936865941571,-0.00628373022770179,-0.0166181189764546,-0.0142750178179645
"1358",0.000530012198390661,-0.0105293773115412,-0.00780370221169358,-0.00688226525108326,0.00693557877540618,0.00262082322879498,0.00424968816603832,-0.00546148757362896,-0.003024769818191,-0.0110518353072266
"1359",0.00196548417766151,-0.00638501249972034,-0.00449446440662193,-0.00506373952748373,-0.00380872206355598,-0.00214705264817849,0.00309262189895554,-0.000866892209536174,-0.00138498223799577,0.000385351197087491
"1360",-0.0032446028501133,-0.00152992714064426,-0.00564329092147065,-0.00482182496808092,0.00374212799667051,0.00289974669267412,-0.00292080523148242,0,0.00838774827586697,0.00346682482868865
"1361",0.0121118133134066,0.00950043211395646,0.0124858047008265,0.0282634587332726,-0.00307972576403659,-0.000839112011936871,0.0136696361555135,0.0138846658243947,-0.0108723413420644,-0.00422251234308701
"1362",-0.0145100203760284,-0.0258045710482447,-0.0134529688978973,-0.0172773908081557,0.0253618780992784,0.00952267599167445,-0.0232782555186061,-0.019971349164595,0.00589325901487858,-0.0185043039401039
"1363",-0.00220094897308976,0.00124665484851771,0.0102274367036133,0.00426228084957136,0.0115743689015806,0.00388448683251652,0.00624590313865525,0.00378454149904472,-0.00190908427597691,-0.00864096828130689
"1364",-0.025176716560534,-0.0211641641090276,-0.0269967956444419,-0.0267904102419453,0.0237402506492876,0.00859022594522219,-0.0253185296304113,-0.0179810911268716,0.0387811976909775,-0.0206023441985491
"1365",-0.000468234856353389,0.00699534906713573,0.0115607243241391,0.00436082671554128,-0.00790137718877082,-0.00576369326216342,-0.00703865994956177,0.00383912265542175,-0.00114281269841265,0.00566352009082416
"1366",0.00757213535192292,0.00315735516891102,0.012571422199571,0.00271360482622907,-0.0133765439889009,-0.00331231379983943,0.0197468052402821,0.00617834589207455,-0.00114421556058042,-0.00362030687199211
"1367",0.0224683825057457,0.0336795302444488,0.0158014348263285,0.0292286479757622,-0.0199842430675442,-0.0065549727509604,0.0213508242923703,0.0362569229353018,0.00044551355762712,0.0185708895967318
"1368",0.000606478564507018,0.00182715746823692,-0.00666645409790068,0.0060478239896391,0.00151919747052265,0.00241638739504979,-0.00486163052442123,-0.00423207961248973,-0.0172381329389546,-0.00673799981177947
"1369",0.0079511908236416,0,-0.00894883640667044,-0.00862513142388122,-0.000239341823295325,0.000741270395980376,0.012538765460409,-0.00510062983160531,0.00148864724919084,0.0031922947283809
"1370",-0.0126968347597149,-0.0112463304647029,-0.004514431924455,-0.0145002646481853,0.00455236999016395,0.00268639987988117,-0.0196208057393861,-0.0150954087703612,0.00407164102815605,-0.0182974890606896
"1371",0.0114906248546072,0.0190595179800142,0.011337667804983,0.0208666691543964,-0.0091432384142075,-0.00535832931201219,0.00935051505101847,0.0118567462956414,0.00708036813156299,0.00486217012124057
"1372",-0.00639509153529139,-0.00904980594131033,-0.00560529915078745,-0.00366888898301065,0.00986947608759658,0.0052944633844243,-0.0047132192540541,-0.00600235162869778,0.00421825367807882,-0.00766118603546284
"1373",0.0106006317050091,0.00700165499973959,0.00789193859509818,0.00710158824788709,-0.00127111044471362,-0.00267846633844326,0.0135531978742438,0.0112133928974325,0.00400970608483031,0.0117837915331112
"1374",0.0102273493394207,0.015719336916173,0.014541144951338,0.0182815637784151,0.00556859116166142,0.00463144054774989,0.00628344194134423,0.012037773223049,0.000570497622820909,-0.00160644505840102
"1375",0.00193791666523246,-0.00922624155559348,0.00220506468815151,0.00205193182157726,0.00537982937767811,-0.000276454587623931,0.00784497589041,0.000855107845812331,0.000570178676385646,0.000804494238004771
"1376",0.00967273578810679,0.0231301895504259,0.00550072210769637,0.0161247127404682,-0.013062673314136,-0.00341331097755837,0.0046637004009864,0.0170991966206899,-0.00487550835261552,0.00844052334810597
"1377",-0.00162119502094915,0.00703782445983969,0.00875270610001855,-0.00327440633044396,0.00494341631579309,-0.00203639848789927,-0.00127633886534662,0.00196109827036373,-0.00757192014324448,-0.0163411536663084
"1378",-0.0224386987772391,-0.0275946994685515,-0.0144547425008654,-0.03662214296607,0.00531582614451409,0.0021332353234631,-0.0156522398117622,-0.0209734768547958,-0.0253253636896495,-0.0214749183216139
"1379",0.00770155613233769,0.011104308152728,0.00666674604021034,0.00318561489911007,-0.0133378980057641,-0.00435002432403864,0.000811058427484745,0.00942637009240888,0.00407837773770869,0.00993788052228783
"1380",-0.0160346805786363,-0.0265405864592144,-0.0154526691049486,-0.0185236860665535,0.0145582487424738,0.00548416677447472,-0.00551234239395271,-0.0116014963177707,0.00733750004807066,0.0102500893865118
"1381",0.00502593799439222,0.00626759954169764,0.0112106946024999,0.00862773029485608,-0.00394235368184015,-0.00221820694731223,0.00440204637809383,0.00973350591015532,-0.00741415216617314,0.00689934024072114
"1382",0.00901664402626356,0.00840873243423768,0.00776080404638591,0.00641541501911869,0.00158315948474463,0.00139002894987117,0.00633003594416137,0.0110574372935379,0.00137601236325557,0.00564301657149979
"1383",-0.00285379004973385,-0.00154418512828847,0.0143014315189569,-0.00478078667732695,0.00244965057354762,0.0032377553875278,0.00838722222409261,0.00168291236512275,-0.0116469212635357,-0.0108217008893704
"1384",0.0249267197852203,0.0423755014122453,0.0206069290425508,0.0443021618512902,-0.0130071964255044,-0.00461092578916078,0.0227123319553453,0.0296750216100696,0.0274081358343303,0.0433548923793641
"1385",0.00301279809010446,0.00919876534153641,-0.0031877741801285,0,0.0103176656727051,0.0046394794984761,0.0106352881113914,0.0103317404693373,-0.000644410069663981,-0.00194172110753565
"1386",0.00659244787266311,0.00793882221363895,0.0127929651842373,0.0199336765143707,-0.0076850106527151,-0.00249371795371234,0.00557089609074812,0.00430574058887601,0.0152815208016381,0.0280155820911756
"1387",-0.00451168615364039,-0.023920534508499,-0.0126313724759237,-0.0105238472602107,0.00510941090223671,0.00268496958397169,-0.00461670828126404,-0.00911037324150166,-0.0113045466840351,0.00378503751243242
"1388",-0.0095035907698483,-0.0128511831857973,-0.00426449343705559,-0.0182324830183368,0.00929386189918868,0.00350935819506581,0.0013914004835649,-0.00432674022920509,-0.0126540730252988,-0.023001542465737
"1389",-0.00125501206677525,-0.000605457782511643,-0.0053534541417688,-0.00361122147411774,0.00881507075726229,0.0027602355655183,0.00200725855901496,-0.000814736796939663,0.00214680882813312,0.0177537984865639
"1390",-0.00871987400918139,-0.00424122988799724,-0.0107641379950102,-0.0111311163610279,0.00202848005724121,0.000459069412934721,-0.0118646509387116,-0.0103289735121278,-0.0122695344448635,-0.0128934580304473
"1391",0.000148995837947696,0.00365092787887789,0.00217637679979665,0.00523545495888911,0.00124574995635185,-0.000917621130921642,0.00155945597414564,0.0107115671484312,0.00552094007969539,0.0111409573662571
"1392",-0.00484500966052104,-0.0103064440822986,-0.0152009977945259,-0.0166663003474388,0.00707572101891207,0.00229569347613023,0.00435932542060646,-0.00625035190354084,-0.00261460871251018,0.00227960414753747
"1393",0.0167774705967902,0.0159266611428115,0.00992306703978874,0.01933255117251,-0.00262480292929945,-0.000824703902611579,0.0108511690730209,0.0150398692909448,0.0101579595034524,0.0121305097542026
"1394",-0.00235717828992599,0.000602940295432841,-0.00436679122467676,-0.00233856700574964,0.00464471033455927,0.00220044395761465,0.00383339025486018,0,0.000454184510537026,0.012359496595415
"1395",0.00686696115568353,0.00421800089917945,-0.00438609955245506,0.0132813861536187,-0.00785977019279493,-0.00256111546961746,0.00840229531483683,0.00942874649218162,-0.00479868988009313,0.00110978658825989
"1396",0.0074073025217285,0.00690084996753426,0.00330384751033819,-0.00257023773101361,0.000543475468058219,0.0010086292875231,-0.00772601617814961,0.00400338786528254,-0.00273667816031353,0.00886924934503464
"1397",0.00262057944025629,0.00953512418596669,0.00768397690326661,0.0092761570199591,-0.00256172622540263,-0.00146591453959155,-0.00839701580605545,0.00318964444954251,0.00215617114362288,0.0120879356194799
"1398",-0.00914823963255318,-0.0242030214719924,-0.0239651066031629,-0.0148073351655478,0.0122192640317702,0.00394538613111828,-0.00338737513294463,-0.0116584364486747,0.00189068320867491,0
"1399",-0.0101125074365602,-0.0229884597734618,-0.0133927303965916,-0.0261724487466513,0.00561275603032452,0.00164524450893366,-0.00602509723040223,-0.0131370545777925,-0.00416476220686868,-0.0209916867428366
"1400",-0.00858630898471979,-0.0145512277169511,-0.00904998703929449,-0.00425764854410915,0.00787522568086341,0.0019158250299014,-0.00404092389067501,-0.00869298540770469,0.00320201923284325,-0.0059150056241617
"1401",0.000223689460796761,0.00691167517381874,0,0.0048104271777154,0.00257880462801907,0.000546254427849613,-0.000156180113736859,0.0112358263140073,0.0140046504949283,0.00743779921520837
"1402",0.0164973474508991,0.0390015708510894,0.0148402192429959,0.0226063011252644,-0.00915571302214235,-0.00309474019790801,0.00811624664666533,0.0181570767953865,0.00706626847904257,0.00184567420582926
"1403",0.0184330476763801,0.0252252776252033,0.0179979538718607,0.0280881767370182,-0.0188616512700311,-0.00721247105319567,0.0113021487163072,0.0159703522140611,0.00491158372363132,0.0103168479898337
"1404",0,0.00029296000004142,-0.00552506263712083,-0.0058182911073178,0.00747198052852016,0.00321873628046898,0.00275576526720323,-0.00314412863171176,-0.000698235399820168,0.00583515216558039
"1405",-0.00699473568058617,-0.00732063806158723,-0.00111111381303985,-0.00458006708058623,0.00200843901134307,0.00174161338041179,-0.00106895535820573,-0.00210221033756652,-0.00597083174614632,-0.0119652153326775
"1406",-0.000871367138367773,0.00147498444217375,-0.0033369860484409,0.00178928831998282,-0.00499875055459398,-0.00364739100200362,-0.00290392363190628,0.00237030402181282,-0.0086267873785294,0.00146794543273732
"1407",-0.00690475238104904,-0.019145963372846,-0.00446439150139233,-0.0117375060234711,0.00566797388586116,0.00239183782326502,0.00107281847400786,-0.00236469896634262,-0.00651021017474662,-0.00842810650609738
"1408",0.0198332806405008,0.044144188571694,0.0112106946024999,0.030983601274621,-0.0161371699507262,-0.0052303402982794,0.00734994658053711,0.0265995366987142,0.00921298873635923,0.0169993723911357
"1409",0.0019374767240885,0.00603960207413556,0.0099778525182852,0.00626124511035298,0.000392152272876256,0.00064570443927936,-0.0028879500232919,-0.00307804324665018,0.00482160067846471,0.00581391130596076
"1410",0.00501378808468966,0.00857630895276373,0.0120748921614975,0.00273746302363032,-0.0128658318363645,-0.00525461974712149,-0.0103656824952605,0.00386010849609764,-0.000127984642457113,0.00758667603917651
"1411",0.00121155167036968,0.000283636420229882,-0.00216941813735039,0.00198532302994892,-0.00532428347601688,-0.00138963619828059,-0.00600767173426675,-0.00589605772402702,0.00127973509905122,0.00286844636302375
"1412",0.000853998136420397,-0.0011336886930603,0.00217413474469863,0.00421137772920765,-0.000719390079334414,-0.000742868913954808,-0.00294450892709708,-0.00567298886288792,0.00325926005263955,0.00822316790061595
"1413",0.00163588563237682,0.000567505563858761,0.00108435455332745,0.0046866767621756,0.00503714401337607,0.00287879716151185,0.00217622298229281,0.00207452551565557,0.00121019169341396,-0.00531922193021361
"1414",-0.000497059977982217,-0.00255177314080857,-0.00216672953267882,-0.00883896778260274,-0.00167059040229778,-0.000648215977063993,-0.000310337825191964,-0.000776561133836062,-0.00757086176992006,-0.00784314027661215
"1415",0.000141986848102293,0.00454814696499239,-0.00108587152639372,-0.000247177652889619,-0.0135468332131135,-0.00491077721491762,-0.000465503098690978,0.000777164649697459,-0.00551317374468951,0.00107795869947758
"1416",0.00113668366987696,-0.00226392002932607,-0.00543467263118924,-0.00148683889733103,-0.0140561331792183,-0.005028961415524,0.00279389587849854,0.000776521205760883,0.00322310309988061,0.00861456835818042
"1417",0.0073784970869275,0.0116279393700942,0.0131148786569537,0.00918088594448818,-0.00852101689860751,-0.00243294558874563,0.0072742749569048,0.00517166083863208,0.0059756664532653,0.00391453712345635
"1418",0.00133820222350933,0.000841076208961011,0.00755101240497846,-0.00491725735522175,0.00487530259185043,0.00121964746438774,-0.000460753970418448,-0.00154349586591818,0.00102199158178307,0.00141799052216385
"1419",0.0000702560614462833,-0.00224080867360832,-0.00214108951566683,-0.000494462837420939,0.00205622574744058,0.000562570549390795,-0.000768668749697721,-0.00206124215967896,0.00344559722150595,0.00460174330616092
"1420",-0.00302433677833602,0.0084221430471747,0,-0.00148332439270071,0.004431312626201,0.000842502345528739,0,0.00180732713605081,0.00998351169984457,0.00916132853008333
"1421",0.000423745745204096,-0.00250528145009443,-0.0010729637947986,0.00049544235359944,0.0165048875678475,0.00776600970121977,-0.000923040707104694,0.00180398707068363,0.0107661712426346,0.00523746664346136
"1422",-0.00817959596772067,-0.00586120548716529,0,-0.00915624866504794,0.00417961955970947,0.00176469193566242,-0.00261786280508214,-0.00565957745595036,0.00840915696314992,-0.00486276892515303
"1423",0.00604272730356858,-0.00364953168185311,-0.00107436051797294,0.000249782030395274,-0.000960241241556803,-0.000463377176117663,0.0038596848777408,0.00129365408939863,0.000494175060190116,-0.00453753155768599
"1424",0.000211774510532114,0.00338101248624145,-0.00322557003784962,-0.0102372521787637,0.00584902193296055,0.00259654548982269,0.00215327433303747,-0.00310098972939921,-0.0037661295069078,-0.00455828677532077
"1425",-0.000988877513745212,0.000561874422693398,-0.00863022342133202,-0.0020179981039008,0.00238954961942706,0.000369992901666283,0.00399009150689977,0.000518592592172018,0.00173523796643993,0.00070453633450196
"1426",0.000777917106895121,-0.0033682576924785,0.00326464251985015,-0.00480298830310555,-0.00437041559865325,-0.000647520299420834,0.000306108123920623,0.00259069966917269,-0.00649593545221427,0.00175991964506861
"1427",-0.00720792929945391,-0.0121090007962444,-0.0184381274536315,-0.0116840831183525,0.00518790532074265,0.00185057559433677,-0.0010698518687009,-0.0108526069303263,-0.000435842840422085,0.0010540966616186
"1428",0.00476860074955576,0.00940715316271978,0.00110484921363141,0.00950910536272609,0.0141333079747012,0.0064635969426432,0.00397733547781898,0.00783666545070827,0.0230500679529013,0.0105300477460186
"1429",-0.000920515965619151,-0.000564976674173767,-0.01324493878931,-0.00560070612875052,-0.00100403065831645,-0.00228755509754086,0.00502810513086249,-0.00596145538963988,0.00158321153584695,0.000347338084005111
"1430",-0.000850535133461228,0.000565296053257835,-0.0123043737124459,-0.00512039764164407,-0.00471256018316402,-0.000368299409963857,-0.000606645664577798,0.00286835909736571,-0.00103354817688583,-0.00486111622344032
"1431",0.0202962544185332,0.0293701448984145,0.0135898732123638,0.0221308049575129,-0.0166510688343403,-0.00681734734233408,0.0078886145726591,0.0176803391220797,0.00352991909841038,-0.000348877680432791
"1432",0.00389515198402957,0.014540521349578,0.0134078235354551,0.0231619816391164,-0.00465415381342427,0.00129852553652232,0.00180633692833498,0.0107308455046315,0.0215295228426802,0.0111692034417417
"1433",-0.00568144619692268,-0.00919435067905772,0,-0.0127949933010922,0.00241855451615991,0.000463384207441964,-0.0064604540811668,-0.01238632517752,-0.00682741027276867,0.00138079096165633
"1434",0.00278738276269208,0.0136462781348325,0.00441015452400273,0.0119638701009683,-0.00627367980351234,-0.00185185895943396,0.0039313163852015,0.0104942239969295,0.00364636873408197,0.00206822407648244
"1435",0.00333537098310832,0.00376970380181785,0.0109770697479616,0.00443341422068144,-0.012464686110171,-0.00491628037736169,0.00376589492732715,0.00531929257058739,0.000119142350892609,0.00515995919531664
"1436",0.0152360386727424,0.016094412699412,0.0162865607119487,0.0269741308403368,-0.00393422587470904,0.0028894433334592,0.0121546816101326,0.0191481166375407,0.0201881850903787,0.00684463933566049
"1437",0.00443486859915843,0.0116156204712452,0.0106838783857475,0.0117000718393163,-0.0265775751124477,-0.00938843933950373,0.00518932839994979,0.00321406405807756,0.00286034093585119,0.0105370807807292
"1438",-0.00339617514406365,-0.00443650048557753,-0.00951385478952216,-0.0108569917863521,0.0120031034843657,0.00206493880511727,-0.00471988668730583,-0.00936428986245597,-0.00814906272149485,-0.02758157108499
"1439",-0.000817745394530833,-0.00786374309444249,0.00213468936497718,0.000477701819248999,0.00501180423220515,0.00252851231467166,-0.00859507820054628,-0.00273631916216699,0.00774652022581646,-0.00726389441688557
"1440",0.000545464433923115,0.00660508191946541,0.00212947624830773,0,0.00656593219721824,0.00233469032377731,-0.00463392925474715,0.000498828683903829,0.000116491962983467,-0.0146341610358031
"1441",0.0000685836597102973,-0.00839885274062646,-0.0106265381702113,-0.00596250558209765,0.00247717130593283,0.000559451085171192,-0.0117134214408509,-0.00299178758538921,-0.0015721671837613,0.005657667601356
"1442",-0.000418308233238962,0.0015880712191374,0.00537033717811597,0.00239910734678106,0.00115311359465897,0.00214187047108583,-0.00030390017314641,-0.00317904418026893,0.00285767771121659,0.0066807125953503
"1443",-0.00150797996072016,-0.00369993486325482,-0.00213675745734909,-0.000957460615984118,0.00781591700216633,0.00223051766602889,-0.0010640776288332,0.000759627789736594,-0.00529195140123473,-0.0104784481678606
"1444",-0.0106422270025381,-0.00822257011552019,0,-0.0148536882210212,0.00987710111272166,0.00370946102862213,-0.014678656648721,-0.00758749537509373,-0.00163694238578882,0.0010589336079363
"1445",-0.00562096167485648,-0.0131049852496923,-0.0107067561267455,-0.00462057108295599,0.0107511686092721,0.00415707666344978,-0.000933860052285018,0.0033131095878276,-0.00562163130241533,-0.00705219856480976
"1446",0.00942131346366937,0.0121949529741814,0.011904885313784,0.0158806603788189,-0.00711755455449592,-0.00211619099076843,0.005453111523952,0.0099058082839476,0.0148989931676462,0.0124289901219379
"1447",-0.00463196864659321,-0.0222220543855541,-0.0192512632910063,-0.00601235160207336,0.000563866654015088,0,-0.00232421094171054,-0.0128269745680026,-0.00261110021146815,0.00596284678055925
"1448",0.00263947658316077,0.00930988484172368,-0.00327151453660168,0.00991988350436013,0.00371082029073877,0.00185603942877921,-0.00714515181224562,0.000764270105686027,0.00232703474505236,0.0013946092478001
"1449",0.00103903754091195,0.00623969635427435,-0.00437637809404023,0.00143779646443165,-0.00136662604652504,-0.000645269061114506,0.00844806553396249,0.00229152648684305,-0.00110271639514203,-0.00522287761086537
"1450",0.00408312411457845,-0.00269611525599012,-0.00439555249921031,-0.00669867256048728,0.000322501064830005,0.00101438855763192,0.00294786876210229,0.00101592058170197,0.00180126664260527,-0.0171508047357199
"1451",0.00716779947889701,0.0121654879774173,0.012141214804759,0.0103563039966383,-0.0124713202767667,-0.00396094776146594,-0.00371244012117378,0.00888086544825351,0.00696013556150743,0.0217237170535389
"1452",0.0000686709217712078,0.00213683644270812,0,0,-0.012953840583724,-0.00453143321798088,0.00434707066300088,-0.000754428372629623,-0.00570247102296839,-0.00522833851815707
"1453",-0.00342127238142054,-0.00799605040824558,-0.00545242090928855,-0.00881997896890641,0.00841888433106019,0.00325095020229571,-0.00417375408050402,-0.00402713050699455,-0.00330200449837803,-0.00280311720481063
"1454",-0.00988756565149251,-0.016388741227483,-0.0164475928327339,-0.00745524928425101,-0.00180058770956759,-0.00203702136738726,-0.00434656428897884,-0.00657061032358741,-0.00616098797743125,0.00737878512213519
"1455",-0.0063801843438015,-0.00273160171134967,-0.00780365151421436,-0.00605774359870104,0.00705200470726619,0.00241278050947269,0.00124745371317925,-0.000254251110860748,-0.000877296892294877,-0.00174399536590708
"1456",0.000558601918921209,0.00986021876935705,0.00561779918982652,0.0092636693723589,0.00692131573844335,0.000925706685973582,0.000155568846274212,0.00610684694241126,0.0028097109063383,0.0115304929006563
"1457",-0.0032783790943085,-0.000271029016738811,0.00111748006150147,-0.0031399186961516,0.0025066693468998,0.0000924646215818559,-0.00435927467731001,0.00126432473700544,-0.00735471018279843,-0.0138169849865292
"1458",0.0083275553047939,0.00922390787120708,0.00669625417139952,0.00581517431082901,-0.00225854741228748,0.000277217673101848,0.00672398962544674,0.0101036412822832,-0.0100552276849962,-0.00490368285955811
"1459",0.010133227990123,0.0185484779269525,0.0144125796813832,0.0103589432053195,-0.0138247279300401,-0.00471470543078023,0.00465998672521284,0.00975234513770418,0.00635575860923931,0.000704040312520915
"1460",0.00453530691387249,0.0102930273380484,0.00546436969159902,0.0078684726895053,-0.00926395431772209,-0.00631619984920284,0.00154602634486478,0.00990585874475691,0.000708269398043582,0.000351663888966014
"1461",-0.00259910339667624,-0.00548587933986799,0.0065217245563165,-0.00283899935475362,-0.00612324431382238,-0.00177569164445024,0.0094162719490305,-0.00662096300178028,-0.00442373499449178,-0.000351540264949435
"1462",-0.0166646527108411,-0.0133964728511849,-0.0129588424284125,-0.0154215464532195,0.0135710205307955,0.00421360817238869,-0.00932843288809782,-0.00987407105480886,-0.0107825823536826,-0.0151249139891453
"1463",0.000139522811618331,0.00559097338366477,0.0142233220973789,0.00963903636023078,-0.00640693459668562,-0.00335680760082646,-0.0035503068602315,0.00772850930456581,0.00365335686857904,-0.00464283041474622
"1464",-0.0138763298470689,-0.0238284447470438,-0.0204963628675494,-0.0205251321860659,0.0143018291078627,0.00477135842357002,-0.010069985004666,-0.0113802785143957,-0.0128297468333961,-0.0121995151716672
"1465",-0.00282867817484711,-0.00135586236275553,0.00220264848086082,0.000974724708432406,-0.00986202292396376,-0.00214159042409345,0.000625900001292035,0.00400418139752623,-0.00344551788743641,-0.00290588105193434
"1466",0.00290773633349772,0.00624674819544091,0.00769229495847013,0.0109540582056566,-0.00510376817413183,-0.00363956590855008,-0.00437885579781316,0.00822516052974898,0.00703629135608219,0.00255005608008707
"1467",-0.000565908707011231,-0.000270086061805341,-0.00545242090928855,-0.00770527649866481,0.0147278308472183,0.00636883973739533,-0.00581233628621547,-0.000494284633097086,-0.000542169605055598,0.00218020271517072
"1468",0,0.00242986728072259,-0.00657902466691707,-0.00145573670700361,0.00587081325823058,0.00409517651553482,0.0112184280703278,0.00766733757462146,0.00542402843348522,-0.000725227892248381
"1469",0.0104707322679849,0.0115807426823988,0.00993373546382004,0.0162818170194967,-0.00818735595197595,-0.00199523553030123,0.00109352876776625,0.0108006098938316,-0.00455550554989503,0.00181427353995822
"1470",-0.00889160612074957,-0.0122471527282717,-0.00765029152251251,-0.00526053866486642,-0.000735859964324792,0.000837050166398123,0.0067114595818154,-0.0111707254471298,-0.0208948085369804,-0.017022771955908
"1471",0.00204833507466806,-0.00377359848341874,0,0.00480775779528875,0.00564343436098369,0.00241544150015027,-0.00744191818189344,-0.000982239660393569,0.00387447710180266,0.00847457402154794
"1472",0.00782531791080365,0.0113637796250023,0.00220264848086082,0.00789485387497679,-0.00943428456984863,-0.00454207449799182,0.00218694557264065,0.00958692930735849,0.0188078605356334,0.0179027562684033
"1473",-0.0226636357496987,-0.0160515259487922,-0.0120879411595032,-0.0163782556023041,0.0181459724137567,0.00838093052686828,-0.00498771012733334,-0.0126613766373163,0.00114252553561278,-0.0186646826118815
"1474",-0.0120241774175222,-0.0108753245626448,-0.00444949388923732,-0.0125482167699508,0.0148387128878156,0.00443241511191861,-0.0101815798529228,-0.00838483182877592,0.00900954985255731,0.0014629624526632
"1475",0.000869283100891627,-0.00329874968404076,0,0.00195496181883659,0.00111256531895831,0.0000915621447843407,-0.00332347424635682,-0.00174079757925893,-0.00101195306232649,0.00803510311144295
"1476",0.000796296361954552,0.00193099533520802,-0.0100558279548175,0.00365874033385016,0.00166694960816316,0.000643438472338387,-0.00158782267865065,0.00024895576675088,-0.00220480267290191,-0.00471015522293972
"1477",-0.00347169735607467,-0.00330342746848522,0.0011286709957572,-0.00899167969889691,0.00332851595508421,0.00119488529052125,-0.00318041593677076,-0.00423397495248545,-0.00209012246205054,-0.00182014263204167
"1478",-0.0134988705050264,-0.00938938219204155,-0.0124013197833592,-0.0154484896636108,0.000947554009210316,0.00027471119653466,-0.0194640617219511,-0.0120058856355381,0.000239335718515754,0.00291761361802267
"1479",-0.00169187717126806,-0.0011151466995617,0.0159818394618183,0.00348677185976443,-0.00197247258003919,-0.000458475516547652,-0.00439310379088376,0.00759494866578736,-0.00628217665598985,-0.00400002006035627
"1480",0.00493739402803306,-0.00558199334762322,0.0179775386394752,0.00297854830426547,-0.000869948573488766,0.000642460691807845,0.0114397443680287,-0.00175873012116268,-0.00126432057954895,0.00438110108307055
"1481",0.0202392346707949,0.0224529541557215,0.0143486314020234,0.0175697757706275,-0.00561814369490243,-0.00201772274577827,0.00937139036459045,0.0148505513167105,0.0119965634194428,0.0189023340870691
"1482",0.000430952795422046,0.00329398000679126,-0.00217619123142432,-0.00194556940982626,-0.0100273502150404,-0.00413569851110573,0.00624304192320624,-0.00248052829848355,-0.00285933171082775,-0.00677854216455243
"1483",0.00186782513159645,0.00355663610067136,0.00109051517737213,-0.00194927464105199,-0.00056238242057749,-0.00147673206055987,-0.000636513747633405,0.00124317722001122,0.00101558636128574,0.00431032299677248
"1484",0.0136250618507676,0.023991332135521,0.0119823520502067,0.0163574608303036,-0.000965383453472413,-0.000554284940603944,0.00811884492630033,0.0144029579269298,0.0122344415401581,0.00357656282013474
"1485",-0.00212230546113634,-0.00213000957780085,0,0,0.0047498215250088,0.00166474351645163,0.00142090720597632,-0.0019584144722552,-0.00106130534130477,-0.0014254239409307
"1486",-0.0051043794881096,-0.00586969355570865,-0.00538211489022744,-0.00840731963180796,0.00392616887995234,0.0023078150291127,-0.00536101399433353,-0.00220755362385805,-0.00424946012952976,-0.00142760560061006
"1487",0.00805227314150825,0.00939338286364833,0.00108246923691024,0.00557160306334792,-0.00143622804029753,0.00128978278707148,-0.00174368567246574,0.0054077049006489,-0.0128030579715404,-0.00321664961115631
"1488",0.00466541418439692,0.0090400041252412,0.0118917974838957,0.00722722995611491,0.000159916972344964,0.00101167036932703,0.00651082575012918,0.00831315541169042,0.00378258774333373,0.00681249553246777
"1489",0.000211187595117845,0.000790545208065874,-0.0032050147206879,-0.000478300940558452,-0.00271742982915513,-0.000183680437103928,0.00394471762304716,0.00193996868700186,-0.00675912218754549,0.000712314306763551
"1490",-0.00492443902698414,0.00368616415509915,-0.00428749934388206,-0.000478615641374303,0.000923573065682248,-0.000396172396354921,0.00282881998800533,0.000484210407111663,0.000481794631464139,0.00249106907856311
"1491",-0.00141359820906717,0.00524683074521715,0.00107655147766761,0.00287266826096522,0.00577525107752397,0.00174913707564728,-0.00125367146795685,0.0021768935461659,-0.0102931857493174,-0.00887467772603245
"1492",0.00176985759033399,0.00182682718128757,0,0.0107423622409479,-0.00047830439338381,0.000827228243152067,-0.0026677224127184,-0.000482703327611578,-0.00182461381613697,-0.00107455759836994
"1493",0.00339200849163834,-0.000260724364321119,0.0053763575596999,0.00755815053337194,0.00215462825920354,0.00055115747276191,0.00881051725061233,-0.000241652858283703,0.00231540952703546,-0.00896381185338879
"1494",0.00302880138430295,-0.00286595971637416,0.00320865534414305,0.00304717821455625,-0.00923638343279098,-0.00284483289653725,0.00405498258866688,0.009420201743217,0.00401218237082057,-0.00108533151390944
"1495",0.000421523219162445,0.00130652500053552,-0.00319839280397993,0.00560883081859753,0.00442014894088993,0.000920634315046742,0,0.000239528732159267,0.00387502412509044,-0.00217317058423616
"1496",0.00680820421126427,0.00887250801570216,-0.00106952138256944,0.00511291838411365,-0.00760133757825043,-0.00193159326763692,0.00124255101095683,0.00310979879466089,-0.000904758729105781,-0.00181478263702284
"1497",0.000487896913103247,0.0043974186261746,0.00428275722714333,0.0030057201057696,-0.011610159202579,-0.00423778130824115,-0.000620462505752206,-0.000715019896269209,0.000724479350117102,0.00472724539946046
"1498",-0.00613204938539036,-0.00283310263868219,-0.00426449343705559,-0.00438004211635146,0.000734502517175217,-0.00194307432243179,-0.00667484827655729,-0.00548936684256296,-0.0084454905363941,-0.00904819863907314
"1499",-0.0037155290256996,0.00490715445341583,0.00535354543584399,0.00439931128506288,0.0074988627809911,0.00222494894913483,-0.00125029305726321,0.00551966631581902,-0.00146005966599916,0.0062089023060381
"1500",0.011752234349905,0.00429216761941187,0.00958456521858886,0.00253572248028466,-0.0149673180652513,-0.00527243147067458,0.00625867712194306,0.00811427190854497,0.00188872838942511,-0.000725868225068038
"1501",0.0111287501177466,0.0087539327082895,0.0150335175673968,0.00698596018352071,-0.010185113158596,-0.00390575974266483,0.0102628364109292,0.00639225808861954,-0.0143517390616426,0.00254264592044251
"1502",-0.00742967624533764,0.000765651235798748,0.0157563365268123,-0.00045922760172179,0.00331903570386149,0.00140009683125175,-0.00140243409231555,-0.00352887400677682,-0.00240621912134487,0.00362325082674775
"1503",0.00575253200524561,0.00586574662165784,0.0134435446151784,0.00597567845776781,0.000165925271376821,0.000652831180996571,0.0113905742891893,0.0144006346534318,-0.0121219987368173,-0.00469318791637974
"1504",-0.00907717100940075,-0.009381078289873,-0.0061223707446586,-0.0114234099110972,0.0109148975184592,0.00270202688321608,-0.00308545756531109,-0.00667216221186828,0.00375637647921812,-0.00181354069069395
"1505",-0.00308111462466332,-0.00204773044143824,0,-0.00208019057927866,-0.00179962474684625,-0.00102233476730262,0.00139240871397672,-0.000486944254985633,0.00180872573057145,-0.00327037887043391
"1506",-0.00421474426343271,0.00102588586509311,-0.00102687331626028,0.00301072935927293,0.00359717740932575,0.00205820710176208,-0.00494499759597933,-0.00097421959741284,0.000996164892173024,0.0102077748250822
"1507",-0.00134044046847726,0.00435564284344436,0.00102792886898695,0.00563557357667022,0.00335554034454955,0.00204462486838008,0.00124255394177997,0.00316869135752151,0.0023635091576284,0
"1508",-0.0108086279911409,-0.014285684179254,-0.00718684290270233,0.00367476352540819,0.00570909465840086,0.00231879219592024,-0.00604944836818067,-0.00753133217874769,-0.00384717662330147,-0.00288700503424477
"1509",0.0169964356607468,0.0170808303000529,0.00827297066451638,0.0148741955574461,-0.0172736890848283,-0.00527457216836857,0.009207439615883,0.0122401185189969,0.00921895517959803,0.00542888193349578
"1510",0.0256302378914401,0.0145038442917329,0.0246156455163848,0.0196168499908786,-0.0133684455040984,-0.00455826197927145,0.0162360745587173,0.0133007474614868,0.00709785194178858,0.00359966281133017
"1511",-0.00225914464224586,-0.0135440896353162,-0.00900911627651435,-0.00707676717696837,-0.0135495721600999,-0.00514018965736374,0,-0.0152746267665644,-0.0120733040641454,-0.00824960277536924
"1512",0.00439128153657387,0.00711924781462714,-0.00404037052929662,0.00200471400793623,0.00390043064119316,0.000469828966023211,0.00608642931012948,-0.00169642692131189,-0.00471460926888234,-0.00433994176907604
"1513",-0.00273253458221423,-0.000757465801935808,-0.00912792692867193,-0.00755715291450232,0.000422032834494157,0.000563373395151334,0.00151246791222359,0.00315602420433403,-0.00629524424962291,0.00181617565745906
"1514",-0.00287704250056386,-0.0020210921069822,-0.0133059443291723,-0.00895866583672023,0.00658517552525373,0.00243969275244393,-0.00196310570202507,-0.0084705299589064,0.00708778178269132,0.00253807371799342
"1515",0.0025416991606606,0.00101260844068318,0.013485380045313,0.00429371114641208,-0.000922602047609078,0.000561599103245713,0.00378254183420901,0.00488155036257365,-0.000435930498703718,-0.00144667207169502
"1516",0.00794962902943808,0.0174508150271855,0.00818826457731969,0.00877588140718699,-0.00277084313015952,-0.00290033879891227,0.00241175840998342,0.00777264581036441,0.00928401117564914,0.00362186399421871
"1517",-0.0000678104770461818,0.0042256574638142,0.00304558917142628,-0.00803028933594141,0.00892422476535248,0.00319002700914739,-0.000150398625717196,-0.00385590536606195,-0.00567970133793549,-0.004330618978589
"1518",-0.000680186003475636,-0.000742808820559659,0.00607311036809843,0.00427228260132084,-0.00275411762135191,-0.00037366545980122,0.00150421248866328,0.00435494747022047,0.00298022479796622,0.00652420086718264
"1519",0.000680648971379094,-0.00346764339495631,-0.00301812615516106,-0.00425410785036762,0.00460229824598613,0.00243245359473954,0.00465551294232558,-0.0019273248145012,0.00631425680450537,-0.00432122496650611
"1520",-0.000136043560842847,-0.00472263440779253,-0.0121091080158734,-0.00089955163457367,0.00208205343897561,0.00130676495411897,-0.00104657522540952,-0.000482663929676108,0.000553617132795337,0.00108497613651792
"1521",0.00645997460890291,0.0107387530727021,0.00408588357814033,0.00562696563076437,-0.00997359256348107,-0.00456768682405961,0.00224447921368642,-0.00217346311735467,0.00430379358021993,0.00433527532181133
"1522",0.00223007724648494,-0.00222355189682655,0.00406914264200653,0.00223783044768089,0.00772295171422921,0.0028092103877364,0.0059716945156989,0.000967933329632853,-0.00159173547872404,0.00647484275670118
"1523",0.00539310569836537,0.000247270921950093,-0.0101316865400342,-0.00156302606429903,0.0019161392603213,0.000840645614014424,0.00504637280372244,-0.00338475763189894,0.00355633094748486,0.00285914600816461
"1524",0.00160938455704152,0.000495225336670346,-0.00818849483376494,-0.00536785957217278,-0.00149661839379556,0.00046692125772041,0.000147610139136445,-0.00388169743873401,-0.00281047843600513,0.00106912297437733
"1525",0.000268022858154193,0.00569177681447641,0.0113519777059186,-0.00359801955464345,-0.00349753328496749,-0.00167892220682309,0.00118112134737336,0.00487092210583073,-0.0109675199021344,-0.000711914167553562
"1526",0.00562225298337737,0.0135335936542564,0.00714292846781883,-0.00338520483137883,-0.0137041634644582,-0.00663352854514665,0.0041292153926884,0.00581665217061511,-0.00477018962669051,-0.00213755737961818
"1527",-0.00119822906823752,-0.00194215383343743,-0.015197714997943,-0.00701998095141121,-0.00364321647489663,-0.00206860364619132,0.0010280096855213,-0.00578301438742579,-0.00224090266694921,-0.000357010471621177
"1528",0.00393129672947445,0.00510818485156017,0.0133745953942388,0.0111745291536771,-0.00552701753323781,-0.00150812414576618,0.00190730950476614,0.00290855799358947,0.0043671597140813,0.00571428109331551
"1529",-0.00391590215613502,-0.00121013697830907,0.0101522874520938,-0.00473609068055525,-0.00170969788415232,0.000566713673081809,-0.00922522571482942,0.00338290742559799,0.00745386025672823,0.0113635906775538
"1530",-0.00246555876918053,-0.00411917179455235,0.00201020348756686,0.00203936968959839,0.00488183140920984,0.000849042767728569,-0.00576417243901295,0.00120478907646571,-0.00610398290765168,-0.000351118811761197
"1531",0.0102875325912246,0.0104623741643046,-0.00300904447931616,0.00655805663826015,-0.0129849125792051,-0.00339737264216311,0.00668945440982038,0.00384862479504333,0.00155086851521458,0.00386373583612265
"1532",-0.0112409240792436,-0.0276908107266806,0.00100590060269456,-0.0132556102003153,0.0128094372395495,0.00577616107443535,-0.00206725265608432,-0.013419725600041,0.00340664608374075,-0.00349897458315218
"1533",0.0100982225544515,0.00693393914140916,-0.0030149802255145,0.00113862914665597,-0.00888739474105593,-0.00357739935152224,-0.00133211371115882,0.00607268905390601,-0.000246870370370411,0.00386237920578703
"1534",0.000728168143909302,-0.00270531339694569,0.0131048301941945,-0.00113733414484907,0.00819086390909107,0.00302363583528442,0.00177815103551193,0.00048253158881284,0.00265492702775694,-0.00139907150236718
"1535",-0.00132309194220814,-0.0120839710540567,0.00298509208314868,-0.00887948982144138,-0.002222844080213,0.000470709379345902,-0.00473275268251838,-0.00627386383840201,-0.0033869265557418,-0.00385290912519543
"1536",0.00556411439299431,0.00848746243536191,-0.00396833289874621,0.00735113229180984,0.00385658419476864,0.000753425438583921,0.00995669302156488,0.0106844638707497,-0.00166824645744557,0.0038678114512305
"1537",-0.000197683718343833,-0.00594089044978063,0.0109561280143196,-0.000455945668591862,-0.000768513574054053,-0.00103491884958751,0.00102997618840317,-0.00336333040697068,-0.0115739921952223,-0.00350257911454177
"1538",0.0016473895855651,0.00821736078564572,-0.00689642657620981,0.00273776206103071,-0.00247797428377694,-0.00103590386019059,0.00587974143004111,0.00168725156398075,0.00118974329097821,0.00175744514794096
"1539",0.000854974330272595,0.00493946495302122,-0.00396833289874621,0.00500569317731192,-0.00813810239977986,-0.00348852575068415,-0.000438235869599013,0.00553566777858783,-0.00525358687381061,0.000350872390607826
"1540",0.000920132979906896,-0.00737302593652867,-0.00996005017583879,-0.000452830683923322,0.00906845980252569,0.00425704373377145,-0.00394745478187142,-0.00526567120131172,-0.00440111277457822,-0.00140306948977265
"1541",-0.00118171024409541,-0.00321849983353539,-0.00301812615516106,-0.0036236947372561,-0.00290983797081379,-0.000942249018857533,0.00117426534534992,-0.00433105995338157,-0.0163562418810391,-0.00421490567380778
"1542",0.00749464136440081,0.0111776155191265,0.0151362857057811,0.00204558953797052,-0.00497881814428858,-0.00160257270299657,0.00689042582220445,0.0113581206640634,-0.00276061256935711,-0.00388012635360513
"1543",-0.0124634966398858,-0.0132649612572994,0.00298209657503756,-0.00884744625494116,0.00301948893055193,0.00217211736321121,-0.00844514491569459,-0.00740754576320146,-0.025043455545697,-0.0113313996413342
"1544",-0.00607898867928336,-0.016430163462183,-0.0118929762012555,-0.0137331916214763,0.00584844679675656,0.00197935526484638,-0.0077825513223222,-0.00698098047563001,0.00779181843909371,-0.0114613456196369
"1545",0.00977286563793056,0.01518636377259,0.0160480397902598,0.00440929989400596,0.000684075786048233,0.00122297337267185,0.00858403558137644,0.0050904061790189,0.00229331680950451,0
"1546",-0.0190270306188242,-0.0309150541592954,-0.0138201116175189,-0.0134008463758896,0.0196532170683561,0.00770369725763786,-0.0168746672165797,-0.0159187325090309,0.00895597170062135,-0.00471015522293972
"1547",0.0068454160282998,0.0069463003187662,0.0190190421800092,0.00562053752054714,-0.00578215870602117,-0.00186465814624015,0.00880579953919725,0.0137254369243522,0.0121809320249042,-0.00182014263204167
"1548",0.0125984140645268,0.0166071379573443,-0.00098237905224452,0.0109453463833085,-0.00295049715627405,-0.000466946265418544,0.00769345827193835,0.010880384005681,-0.0105619894343746,-0.00619988201925725
"1549",-0.00197519780302557,-0.00276477852909407,0.00393310377923695,-0.00460739481216654,0.0018599109766424,0.0014020012406557,0.000146902335386168,-0.000717626807934857,-0.0101572551523531,-0.00440368522061918
"1550",0.00329838815725259,-0.00453614681267556,0.00979409998635572,0.00231456676057351,0.00544578501731374,0.00249431927573829,0.00190837042903302,0.00694108961636952,-0.00366011764705887,-0.0070032599178137
"1551",0.00532499831852018,0.004050338697005,0.00581949085816791,-0.00946678405590795,-0.00529820830352001,-0.00233006437243188,0.00747238014051788,0.00499150307261731,-0.000918387550270405,-0.00371197812652269
"1552",0.00895892931578501,0.0115986365884779,0.001928787554907,0.0121212550819274,-0.00287499004679681,-0.00102723941408334,0.00770829621688418,0.00402068631077457,0.000525292176126957,0.00931452061308158
"1553",0.0013614689487369,0,0.0125121316852825,0.00483644100055747,-0.00907328298461429,-0.00317968560234327,-0.00375258192721084,0.00235574846562692,0.00557810061759745,-0.00553713659489818
"1554",0.00181240255111437,0.00672978553609327,-0.0095057852893401,0.00275031240741375,-0.00770117336195753,-0.00384609444721129,-0.00362152057692722,0.00164544590040894,-0.00352407501204921,0.0066815377053342
"1555",0.00426362213777498,-0.000742528101790874,0.00479838477461825,0.00868591916671657,-0.0104350695449205,-0.00508526278084409,0.000581399326773369,-0.00351945766585926,0.000131017091741237,0.0029498120940703
"1556",0.00379559448729117,0.0032210154893384,0.00573069319439501,-0.00543851656911487,0.000958488509732014,0.00047369992204005,0.00392328698316757,-0.0014128106571677,0.00183352751728982,0.000735284073664522
"1557",-0.00224320110666187,-0.00271657897768018,-0.0104462988914017,-0.0113923122887684,0.00722650033842642,0.00274333657283266,-0.00361845315907006,-0.00589492394392244,0.00784363004628963,0.00220426929571249
"1558",0.00141326500604744,-0.00247667696151066,0.00575816427873677,-0.00944900376669611,-0.00103723269163458,-0.000849573534621451,0.000290786196696091,-0.00047416694489355,-0.00343730457957969,-0.00513193244750831
"1559",0.00532383146457804,0.0139029002372384,0.00572530497864476,0.00418801113512202,-0.00302822286653992,0.000284079262128811,0.00537307849412838,0.0163741704167963,0.000130085900557519,0.00736920964057641
"1560",-0.00132012355340672,-0.00171412828433348,0.00948774738854241,-0.00903625848257017,0.00468630104199663,0.00349282267741358,0.000433384126550251,0.000280840070292943,0.00208229447277497,0.00219455661418477
"1561",-0.00551909789573202,-0.0139809254864685,-0.0046993805366824,-0.0112227638029533,0.00760234763159207,0.00329227451929937,-0.00274319748773111,-0.00726501873241892,0.0089610714285715,-0.00583944890513199
"1562",-0.0023231560200726,-0.00248779811604993,0.00566572877348515,-0.00709380124385051,0.00677272843548526,0.0030942725323504,-0.00709437167330351,-0.00613815343068014,0.00450506485696156,-0.0073420437609536
"1563",0.00698581738790138,0.00573602826754893,0.00751159589695227,0.00571534859510292,-0.0111555598341958,-0.00383259395150026,0.00583244975288011,0.00356324858527546,-0.00454899404729647,0.00702653066856218
"1564",-0.00854266646802415,-0.0116541121777122,0,-0.010182189073325,0.00964498551951198,0.00262722353292943,-0.00333418242757877,-0.00591715257645398,0.00566393144313371,-0.0044069196129316
"1565",0.00803298481647641,0.0102863529922406,0.00372804521560588,0.00382793111463187,0.000768059214765637,0.000374604496592434,0.0061089613851677,0.0128571299408773,-0.00447998080000001,0.00184431274578434
"1566",-0.00417739980881782,-0.015644833162757,-0.00928515686388209,-0.00095355996238311,-0.000937804771031669,0.000748074585845249,-0.000670374121873429,-0.00188037942732977,-0.00199291542283031,0.000736442796368086
"1567",0.00800285768212361,0.00479359074485353,0.0093721790162038,0.0143132544650799,0.00119442743850473,0.00102867742621671,0.00744066321120074,0.00894937150634223,-0.00334967781017526,0.00919792752690629
"1568",0,-0.0100431287611256,0.00464216067795009,0.00376283190913873,0.00852078138730361,0.00429598944099219,0.00159329449402823,0.00396803843639804,0.00413650462683246,0.00510390617331535
"1569",0.0030731937303905,0.0071012893135658,-0.0018481802828475,0.00210865494266432,-0.00506972590985355,-0.00185997273864846,0.00462681669119513,0,-0.00585738925169044,-0.00943056091566707
"1570",-0.00395738289226966,-0.00528815239017455,-0.038888779243765,-0.0107552215504261,0.00753196939514433,0.00265888786977775,0.0031663713119181,-0.0179021495649229,0.00142441569616869,0
"1571",0.0049345695519869,0.0108859764552613,0.0125238861399584,0.000472962351652173,-0.00405450372366145,-0.00195415177468372,0.0025825698483315,0.0187024499167037,-0.0144824790131568,-0.00476013385914431
"1572",-0.0101395206780546,-0.00500873900852905,-0.00380589509597462,-0.011811958629437,0.008989806876746,0.00419519996451556,-0.00529488854891025,-0.00720447416718939,-0.0111526410684805,-0.0169242426921778
"1573",0.00405863807020213,0,0.0410696993155999,-0.00286897378981676,0.0119356748144397,0.00399209245962306,0.0146739295337777,0.0203653572296267,-0.00291914689628192,-0.0011226621444842
"1574",-0.00449135656683841,-0.00604057318922213,0.00550469749665328,-0.00239760496388841,0.0201847063469869,0.00314336219367006,0.00269391416430032,0.0142235006692617,0.01676761672349,-0.000749411160418934
"1575",0.00676747855542925,0.000759545532936778,0.0100363757203425,0.00168244560114439,-0.00765356288085017,-0.00322617094097,0.00933257789204278,0.0022620012803205,-0.00425360911267092,0.00299958406858414
"1576",0.0034567950435298,0.00556676552299651,-0.00813010463765773,0.00983689328888548,-0.002461551280175,0.000369870562480168,0.000420607361264036,-0.00112856390036864,0.00775494196227822,0.00635520752959895
"1577",0.0122489855201553,0.0158528881611217,0.0209472515331008,0.00950343887021465,-0.0137357158460055,-0.00415949468432986,0.00588153493749255,0.00610027591895923,-0.0168905443299999,-0.00222887210996559
"1578",0.00327692802070967,0.00569729230253468,0.0115968826104957,0.000941386191936511,0.00191774815052459,0.00111390938155309,0.00487243607464083,0.00381744297698261,0.00199006965174142,-0.00409532978060922
"1579",-0.00245003241830755,-0.000985204270340767,0.00176343077920471,-0.0152834106051503,0.0148998501958413,0.00556322146876753,0.00581899507645955,0.0123046167552618,-0.0470043419992517,-0.0123363959983461
"1580",-0.0231737166186198,-0.0219428139594186,-0.00792238542591994,-0.024355437924744,0.00869311562589625,0.00221319858408831,-0.024931510316102,-0.0227625116244619,-0.087808261642409,-0.0299015704037351
"1581",0.0147629655102888,0.0143686652064248,0.00976048387080675,0.020558360936201,-0.00821170302185437,-0.00285207549647704,0.0158217456790171,0.0174127789445471,0.0113472319145111,0.0105344659073492
"1582",-0.0146112709310987,-0.028081820044775,-0.00702981947953751,-0.0158274372783512,0.0066405641673335,0.00184509705258407,-0.0120986401040037,-0.0111135013193092,0.000527048180864798,-0.0146718133830123
"1583",-0.00625400057522119,-0.000766637782530499,-0.00707961258809475,0,0.00244278517895502,0.000552472491850198,0,0.000449210375425002,0.0107624599519254,0.0105799947329301
"1584",0.00869321585127247,0.00690881314076086,0.0106951237725259,0.0146200760886059,-0.00211152790102631,-0.000552167434531681,0.0115429401741007,0.0146036357877208,0.00871182407940818,-0.00232653110253789
"1585",0.00443835203820164,0.00482847193339753,-0.000881789781316256,0.00480269905559227,0.000732039494237835,0.000552472491850198,0.00139152774479268,-0.00221415799482649,0.0179374989448771,0.00310924862864859
"1586",0.0103088779982097,0.017197942744055,0.00970839714329919,0.00478028281610521,-0.00349760883605277,-0.000644368797508288,0.00583678518167163,0.00199683559687358,-0.00739658480333205,-0.00619922233375714
"1587",0.0006340265114535,0.00795600419465314,0.00611906620306546,0.00594666416657952,0.00253038798804539,0.000460666464185966,0.00317756385269474,0.00442998009871576,0.0108853736526382,0.0109162716021534
"1588",0.00405372985925467,0.00518025498409425,0.00521313376861876,0.00898556209712242,-0.0043157246871095,-0.00110486737847271,-0.00123988077149628,0.00308700868005385,0.0235600933569451,0.0131122044342977
"1589",-0.00176657232757738,0.00294473245117688,-0.00259300036456445,-0.010077302712165,0.00916014048874669,0.0035946764365864,-0.00455009406480489,-0.00395653404562146,-0.00508367559543632,-0.00570989639238018
"1590",0.00669872530499105,0.0149252899403758,0.00606547866943163,0.0104166490903097,-0.00364733640152315,-0.000367725539134112,0.00775716834121454,0.0134626855133348,0.00986444511065376,0.0133996281898012
"1591",0.00238534418669611,0.000482211844776481,0.00775213099799288,0.0142926131058905,0.000569470157083973,-0.000183252047499027,0.00975928734811449,0.0041376211709907,0.00330288819459823,-0.00755569810693069
"1592",-0.00876725416296442,-0.00578299910764435,-0.0111108408593378,-0.0108570722342627,0.0102732338216593,0.00326583218855347,-0.00680629781094833,-0.00303660408589379,-0.011627113213501,-0.0178911993642445
"1593",0.00928761528574618,0.0048471922043265,0.00432137562279733,0.00794012861010418,-0.00129069533170034,0,0.00383737876293466,0.00478567542277286,0.00574018137807242,0.0127906433562244
"1594",0.0101401197795117,0.0125421059562687,0.0137692740736874,0.00834089703470808,-0.0235767116829566,-0.0085285089206526,0.000819435186111939,0.00974281663439869,0.00119784387257416,0.0110984797220384
"1595",0.00254087142164416,-0.00214381012246911,-0.00424450730057169,0.00137878225145793,-0.00248112174872761,-0.0012945659563387,0.00395651964441046,-0.00171536286996199,0.000422253513188808,0.00113548788016282
"1596",0.00506886351284797,0.00429692147835636,0.0017049680565111,0.0071134091459879,-0.00389601560482356,-0.0013889685693157,0.00584321780613961,-0.00536937753405287,-0.0124515587387221,-0.00340260002939397
"1597",0.00455074489770468,0.0125982432598606,0.00851080908052881,0.00774685355119953,0.00158115119068714,0.00120534307459153,0.00243170121731207,0.00539836338513355,0.0148169392072608,0.00455228966012333
"1598",-0.00281579315381664,-0.0103289228880789,-0.0075950522349828,-0.00723508485192481,-0.00257559364950977,-0.000184768327137319,-0.00512116220124648,-0.0124567820546512,-0.0115822611183781,-0.00037763835250948
"1599",0.00325394766463338,0.0040324836070782,0,-0.00774300013526308,-0.0107465911002996,-0.00565177865734601,0.000270729481269605,-0.00282781444177671,-0.00859308299968875,-0.00453344997004712
"1600",0.000795114357152515,-0.00496087251411936,0.0127552258078738,-0.00918097603028245,-0.0076630160817186,-0.00177015976518824,0.00148981197328779,-0.00937789806597511,-0.00838118158820145,-0.00455409573522136
"1601",0.0103340328422179,0.0018993900674098,0.00671691839950772,0.00463300993645577,-0.0108623981256242,-0.00401365082672545,0.00527401402303451,-0.00440335265544656,-0.00447876205556108,-0.00343117818564065
"1602",0.00538635618844574,0.00402797741758065,0.00917446039014802,0.000230619182925329,0.00669179953758792,0.00262432557061643,0.008877909666271,-0.00309617408686491,-0.0230751980708975,-0.00229530155362823
"1603",-0.0046952155566804,-0.00330407768793795,-0.0148760730071297,-0.00345780557129627,0.0103973072002774,0.00476669884739378,-0.00319972613469244,-0.00155291133880264,-0.00401105979309735,-0.00115036996924256
"1604",0.00967686900149478,0.00710391690735346,0.0159396905697937,0.00439504776678068,-0.0126516291479029,-0.00539522976009021,0.00628661549951492,0.0135526159175514,-0.0225221052284915,0.0049904142640429
"1605",-0.0000597926556656914,0.00352733037236264,0.00660589326905026,0.00253347938080717,-0.00119582153230446,-0.000748148021375461,-0.000531574984944938,0.00548007766011782,0.0308994261364461,0.00649353610594772
"1606",0.00143784308697747,0.00234265260103372,0.00574258453074528,-0.00206769783127625,0.00786836264067925,0.00262030062241503,0.00465464968318607,-0.00893846216642336,-0.0165777833251103,-0.00569256107987448
"1607",-0.00741753984765914,-0.00864886427936284,-0.0106037651209292,-0.0110497779943041,-0.0148507372493694,-0.0079350853444754,-0.0247551991284582,-0.0217772157062301,-0.00707407408661687,-0.00458016862487476
"1608",-0.00289301638945449,-0.00495139684092605,-0.042044375095511,-0.00744866985431247,0.00473819121258479,0.00103525491066203,-0.0139811807148518,-0.0179897836236305,0.0202364632372829,0.00460124309412979
"1609",-0.000845860028275247,-0.000710887590332443,-0.018072128359734,-0.00867735019960236,0.00137145100899105,0.000376260012306506,-0.00385441126134556,-0.0137392650922583,-0.00631458282211894,-0.00381682028174757
"1610",0.00598856974372453,0.00497954540165702,-0.00613515197107095,0.00544143168415046,-0.0253425227898287,-0.0117463724369592,-0.00995045765861791,0.00371458225527932,-0.00201846598454203,0.00919547400448573
"1611",-0.00649432900818581,-0.00542708003955095,-0.016754749762145,-0.0127059592322268,0.011243740964908,0.00408891070862549,-0.0199606121748089,-0.0168860293072748,0.0100381822594133,-0.00645409096761351
"1612",0.00369207128021931,0.00711742947932059,-0.00538147427927016,0,-0.00243210492311663,0.0000944979063257634,-0.00954297335363885,-0.0115297565998537,0.013869279628135,0
"1613",-0.014352129011403,-0.0209658219886766,-0.0225425622924923,-0.0181124302767844,-0.00339617467198305,-0.00274581040129862,-0.0122233547909689,-0.0211854185067967,-0.0203364964228931,-0.0118455806241523
"1614",0.00550641128811113,0.0098653198034615,-0.0119926374196364,0.0148059193807522,0.00529903448443081,0.00144542767891109,0.00247520458017347,0.00437747552266643,0.0193398823079434,0.0123741931688792
"1615",-0.00480706067953685,-0.00381226798317003,0.0289449479727573,-0.0121984873150671,-0.00923529999497752,-0.00256360232919961,-0.011617984134907,0.00750615534345589,-0.0093765954646764,0.0038197756843481
"1616",-0.0140008419839236,-0.015067895748377,-0.0381126148910088,-0.0179175851770196,0.0138060462343153,0.0048542386090662,-0.0107257312059206,-0.0206682136922014,0.00214455378672063,-0.00456618679793841
"1617",0.00905330221117606,0.00801324040329154,-0.000943348700596758,0.00838287619647637,-0.000606750657995647,0.00123165624704358,0.0187137977098337,0.00490816409944661,0.0074527373833313,0.00382265631848155
"1618",0.012720418267125,0.00939530976303948,0.0387157823064981,-0.00513466381358507,-0.0178792440944269,-0.007757732134133,-0.000583383077603972,0.0144074614222613,-0.0238042922713271,0.00228477333300514
"1619",0,-0.00167037565841899,0.0127271420735426,-0.0135167034873651,-0.00477196320150364,-0.0024791775713281,-0.00875266337797342,-0.0122769409982993,0.00495200333847534,-0.00379945755776012
"1620",-0.0103158069434524,-0.00980187943890276,-0.0197485687098893,-0.0189335834254751,0.0118983519363134,0.00248533916845162,-0.0153051472997449,-0.0216916755394456,-0.00515157525531462,-0.00877181068797406
"1621",-0.00827696419063961,-0.00120697375777956,0.00274734605917448,-0.00685625312335136,-0.014303127940954,-0.00448135432507057,-0.0146464749327911,-0.00747345314050207,0.00750469043151969,0.00115427429577508
"1622",0.0152085296591704,0.0120859266167532,0.023744094978948,0.0212220533022007,0.015668111419642,0.00756666844075848,0.0304868498108826,0.0256020774277721,-0.00379884543761644,0.00653342551185299
"1623",-0.00627260729558055,-0.00740382688601815,-0.0312219324508749,-0.0157736779082763,-0.00236664837894518,0.0013302025124895,0.00250202059562699,0.00244731375173735,0.00515917432484025,0.00420005822399827
"1624",0.00772169588285476,0.0098653198034615,0.0267034972194538,0.00915767884475271,-0.00527167132628292,-0.00237299499707311,0.00132111806783786,0.00366206223651622,-0.00490953681742734,0.00228141593051934
"1625",0.00790577381936219,0.00333568602183898,0.0170402549700512,0.00428559361115988,0.000530173910610499,-0.000571182711978535,0.00161338583880144,0.00997306468299319,-0.0122598411524305,0.00189678735838483
"1626",-0.0138169021771655,-0.0189979389328565,-0.0123457264638503,-0.0308735033383944,-0.0103282827592026,-0.0137105769950312,-0.0300103492930053,-0.0236025300491807,-0.0116552557460359,0.00151455709395831
"1627",-0.0247782596879365,-0.0326797017266263,-0.0410715202575598,-0.0448072161603192,-0.0164125931457921,-0.00453699590077705,-0.0390886388578154,-0.0434139388238095,-0.0535262900230122,-0.0325141227318189
"1628",0.00321021837811553,-0.00900913007123583,0.0363128574263394,0.0143711343951767,-0.0169586070856812,-0.0105702836844291,0.0117795468947952,0.00489204857795089,0.0117314322286639,-0.00625247726745759
"1629",-0.0126359320570326,-0.015404020121882,-0.0278527920060372,-0.0203152649438685,0.00415144212600027,-0.00245006892792621,-0.00636446103560206,-0.0190053490590819,-0.00895644120856198,-0.00432562145749138
"1630",0.00961389642777144,0.0118642692261464,0.0129392631313476,0.0212823422289956,-0.00891161617000824,-0.00117857826564227,0.0184347972820309,0.0177812040804006,-0.00371176470588241,0.000789878627295737
"1631",0.00990153010961015,0.00726340667183778,-0.00456199362870069,0.0157624394131026,0.00648928874315424,0.00403250294267776,0.0149571863549851,0.010430091339747,-0.0420345181660766,-0.00276239324015415
"1632",0.00586945140412287,0.00463532243386999,0.0245786912884702,0.0200657177367904,0.0102227768115921,0.00538892501944366,0.0178490010335584,0.0198712071210956,-0.0197835392271182,-0.000395720742039196
"1633",-0.00409719328436464,-0.00666489378445723,0.00808638301561215,0.00574703859849124,0.00683719086485723,-0.00116995100406847,-0.00434669922595188,0.00961555232948785,0.0273417193834444,-0.00514652842086805
"1634",0.00585998061648318,0.0118708118577953,0.0124775147653167,0.00311723718968526,0.0020148060623062,0.0003812419186211,-0.0052683269802285,-0.00451131991465659,0.0169590796997812,0.00636692819458662
"1635",-0.000929744692862444,-0.0104563940575166,0.00704224918187535,-0.0178665846074333,-0.000633789819923569,0.000390433821467306,0.0116522091583944,0.00881172522619345,-0.00891599130477971,0.00395407799903147
"1636",0.000433686547834711,0.00128881833931183,0.00087425689020959,-0.00922748670306162,-0.00299134365911535,-0.00195242806885287,-0.00433816837906853,-0.00349394605683417,0.00574756337157267,0.00905876382185755
"1637",0.0107890442463097,0.00180182171182897,0.013100564499984,-0.00638647598861242,-0.034087578933868,-0.0168228450358633,-0.0105166867412206,0.00776346752412627,-0.0219480043390426,-0.00234196863799574
"1638",0.00570473799690929,0.0107911402618202,-0.00689654573150222,0.00133902327163682,0.00969303207696148,0.00586992684413201,0.00394750913589315,-0.00422447443570417,0.0120247781192235,0.00508608309389769
"1639",0.00719719411958519,0.00279616327561527,0.00520816472001218,0.0131050621990056,0.00102563261884203,0.00168095100710208,0.0127044353975891,0.00798598209222812,0.00928793390866134,0.0062280993616175
"1640",0.000363471968898743,0.00709751656211721,-0.00345419272253633,-0.00950353716479868,-0.00782146296575814,-0.00355432813612544,0,-0.00594209620844754,0.00273581488801655,0.00309481492883301
"1641",0.0136207322027393,0.0279388484478029,0.029462661729603,0.0490404279067358,0.0117307108325624,0.0100079054249544,0.0276284955982817,0.0328767427994021,0.0272013318032576,0.00501346891729848
"1642",0.000417868417277534,-0.00759086526658115,-0.00168330611568546,-0.0106709150703924,-0.000834656768354702,-0.000785245940304713,-0.00653956457946947,-0.00795752326318011,-0.000885391192617324,0.00383732509349644
"1643",0.0038211472219285,0.00444150241394259,0.00927470317361445,0.0102722472669285,0.00529129383064975,0.00314189506376494,0.0036565583918351,0.00607677540435358,0.000402827690393126,-0.00267588302880972
"1644",-0.00374702836924989,0.00122798975427418,-0.00835409024024891,0.00406722177253416,0.00341683613332089,0.000489484039752908,-0.00160284803754096,-0.0026578324566997,0.00571749879207606,0.00114992905154732
"1645",0.00256707565524139,0.00147226647840215,0.00926705508514059,0.00911424638519232,0.00184075099186143,0.00440217800733622,0.00525538882883247,-0.00314906988418795,-0.0125710546286417,-0.000765765091293669
"1646",0.00547752618809327,0.00857411242642114,0.00500825547660644,-0.0117914841510125,-0.0124931135965726,-0.00467511258834841,0.00624461401564358,0.00267326363411158,0.00559521569899446,0.00421458075059888
"1647",0.00177638353548404,0.00291473354224503,-0.00747517932105102,-0.00279257380989151,0.0158133924190658,0.0054798928842823,-0.00101044727156308,0.000969198458304676,0.00887024419207738,0.000763017835870849
"1648",0.00195099227917428,0.004843820304264,0.00251064902485565,0.00992874603158334,0.00146569387068451,-0.0000965098518954655,0.00288918862425547,0.00508479973127218,0.0298137236846479,-0.000762436083540319
"1649",-0.00212366996856916,0.00168711319609227,-0.000834849474449895,0.0108393119972805,-0.00420615433241645,-0.00116819623092712,-0.00043192452522367,0.000481785201643214,0.00675264690321775,0.00152611420787818
"1650",-0.00366575577239758,0.00288746995425315,-0.00835409024024891,-0.0102241788593602,-0.0126725909193552,-0.00672405215228167,-0.0194552227242437,-0.00866858387867486,-0.0171922278903276,-0.00799996926074609
"1651",0.00243273048331227,0.00575813688818094,-0.0185342045221828,0.00579461898864708,-0.000372277428990153,0.00147114246818481,-0.00117588003676494,0.00364352898287068,0.0093347581737977,-0.00115205797759044
"1652",0.00106546936756202,-0.00238567252052324,-0.0231760235723585,-0.0022543758052338,0.00614051106584013,0.000881742326349189,0.00264874818265137,-0.000968036199426758,0.000854907917228864,-0.00615151468866593
"1653",-0.00307473439632211,-0.00382585900137467,-0.0219683597810465,-0.0125532788359511,-0.00730478811915958,-0.00205525257778005,-0.00792484780178826,-0.00823647325457566,-0.00240719057623229,-0.000386841912370151
"1654",0,-0.00336057510611454,0.00898499020842425,-0.00228828326764086,-0.000372945362871246,-0.000294004482731425,-0.00118363078164296,-0.00610635735291465,-0.00272441813089119,-0.0034830042132139
"1655",0.000712127664696638,0.00602125766980777,-0.000890605114578058,-0.00586139992940049,0.00363474597781699,0.000686584262123979,-0.0137736964865748,-0.00442366176214148,-0.00124879805060862,0.00699035586535879
"1656",0.0115579525150651,0.0100549116264639,0.0276292265278906,0.0182001467625308,-0.0192685861842244,-0.0088256657572644,-0.00555645423692896,0.0118490250204111,-0.0105501563812922,0.00231393010372782
"1657",0.00169925100091928,0.00568876493276882,0.0156115753733674,-0.000251675326431222,0.0110099390708427,0.00851824257187306,-0.00437922324031026,0.00146340913089182,-0.00197456755410652,-0.00384769978730604
"1658",-0.00146206636767032,-0.00259276043129408,0.00256174611522697,-0.00629526815720616,-0.00769811374149587,-0.00314293796815335,-0.000606676622038282,0.000487289719014239,-0.00522320350408989,-0.00502117525665891
"1659",-0.00568282713786983,-0.00165402516931989,0.000851725497169165,-0.0126714283417891,0.00293293136328243,0.000295708739757927,-0.00349058791389867,-0.00146098121737848,-0.0137628961120818,-0.00815226196392715
"1660",-0.0032401628163653,0.00142057683530816,-0.0187233016796093,-0.0107803827783882,0.00745255945564183,0.00364389392712727,-0.00411228608999747,-0.00658355891554208,0.00145197223963889,-0.00665361032499945
"1661",0.00366458102524336,0.0103992973707108,-0.0052038179852143,0.0192010395684115,0.00271489915053547,0.00147201932894525,0.000917791143417057,0.0112910272634863,0.0218284249403395,0.0051221547324638
"1662",-0.00288556272653429,0.0016370728904409,0.000871945672805019,0.0020365824278894,0.00158750775390559,0.000685863674928955,0.00947261062368465,-0.00169863795738878,0,0.00705608126312685
"1663",-0.0011817360889117,-0.00373642619948444,-0.000871186045901973,0.00940064180033429,-0.006806188960777,-0.00195816464970011,-0.00817299955347028,-0.00705125135301332,0.0178937725217267,0.0120669074580908
"1664",0.00295688726639209,0.00609461460704042,0.00871843148397633,0.00604048555133629,-0.0144558710981335,-0.00902706788324559,-0.013734026756545,0.0017142128824168,-0.0107643998000311,-0.000384530976713426
"1665",-0.00512963218369056,0.000233271051729211,-0.00518592388217209,0.00325248841265435,0.00152456510604515,0.000891234193523438,-0.00216634248442293,-0.000978020277415448,0.00986380162617517,0.00807999927135161
"1666",-0.0139857786553237,-0.00512486891178765,-0.0139008237061168,-0.0114713907898357,-0.0135046931083616,-0.00553939038041251,-0.0189175998456204,-0.009052724211431,0.0208527286821705,0.0095419721382568
"1667",-0.00330572214294322,0.00210709890530003,0,-0.00857712870188931,-0.00347115923280239,-0.00388027844643979,-0.0230759486043257,-0.000740967597493425,0.00675829589553811,0.000378066669932675
"1668",-0.00639203872979721,-0.00887829510489568,-0.00264319723553175,-0.0188296001810091,-0.00870635500879102,-0.00429339967699049,-0.0135897402391688,-0.0113667498775476,-0.00429934372757068,-0.00113377136863213
"1669",0.00491604523448363,0.00353583951846947,-0.0088339580078437,-0.00181505972626828,0.00770976359493414,0.0054160342000138,0.0234540846649962,0.00324931768012826,0.00333309610382138,-0.00189184165773648
"1670",-0.00616031944190476,-0.0112753951159013,-0.0142602379000465,-0.0233827719262226,-0.0109431152847898,-0.00628458845473312,-0.0020833652540776,-0.017438695237214,-0.00286893173731062,-0.0011372096858524
"1671",0.00911539438369591,0.0125920562628712,0.00632897260596121,0.0162275350821492,0.0101825397867965,-0.000401477195545841,0.00562068281018702,0.000506668509453023,0.00560302082818853,0.000379579586898826
"1672",0.00337188497697238,0.00610056452878127,0.0170711468175881,0.0117802683819461,0.0108559273515014,0.00562294974355337,0.011657635051729,0.00734952830959124,0.0157367369284953,0.00796658499444414
"1673",-0.00372088640207113,-0.0062967481732854,-0.0114841602506172,-0.0108667565212036,0.0049860892979301,0.00199775413672709,-0.00378822226332498,-0.00654084946190403,0.00407711656384513,0.00564542635091381
"1674",-0.0160839620001292,-0.0194789631457647,-0.0107238646146997,-0.023018554706848,0.0125937544563368,0.00568079046222492,-0.00301108279074047,-0.015700085371021,0.00959765986558136,0.00973052179638567
"1675",0.00355113377052851,-0.00215423583878083,0.0027101292988978,0.0021417880112673,-0.00810295423610408,-0.00406296950517115,-0.00476776532194156,0.000771668135262527,-0.000292453382084168,0.00148263579272623
"1676",0.00158598342264682,-0.00263834253461592,-0.000901136577268646,0.00801513476364302,0.00797964466462919,0.000995081334079329,0.0015969874473758,-0.00128518378685394,-0.00614448070359619,-0.0103626668671772
"1677",-0.00316758596865285,-0.010822811208879,-0.0198375839784912,0.0076858944337288,-0.00113055488793756,-0.00188888114059627,-0.00765294477654577,0.000514772241088313,-0.0091999708986521,-0.00299180861046588
"1678",0.00452182610058549,0.0143452251368408,0.0248391710112228,0.00631253669967435,-0.0141049529216724,-0.00567526432388799,-0.00835484044470325,0.0128635025918509,0.0133709929197368,0.00525124106240105
"1679",0.00827304325866596,0.00479374861408721,0.0152602179547852,0.0177729938897557,-0.00220607798538097,-0.00331033495665567,0.00712900801496064,0.00457172096021208,-0.0129012903225523,-0.00858201128343494
"1680",0.00126702284693714,0.0004768252372922,-0.0026526198368314,0.011813088873446,-0.0139441051024549,-0.00764894744197475,-0.00852654590125845,-0.00176975985197381,-0.0182682825406718,-0.00225815504595728
"1681",0.00048205893524389,0.00643808257891942,0.00354623325779424,0.014720932620836,0.00497358511320356,0.006085603315787,0.0183352922539344,0.0032928637354348,0.0147503558566646,0.00565820345158907
"1682",0.00957620300279172,0.0106608122695004,0.0256182259356033,0.0262632022489044,0.000485223522156186,0.00201568284421394,0.0197578335547435,0.0217115544546453,-0.00178896765362513,-0.00637662282010609
"1683",0.00739682084720683,0.0128926767204001,0.0077519656527163,0.00755532090131994,-0.00698335172209175,-0.0046273785296852,-0.00124996388395848,0.0113662142541457,-0.0162049057962839,-0.00906001565387571
"1684",0.00313864968205291,0.00740537510213168,-0.00683741036035046,0.000725864000943321,0.00888824425778578,0.0050535846890285,0.00688372383536406,0.00464233047708573,-0.000303689073034463,0.00152390635694055
"1685",-0.00265634083385258,-0.00413506630123683,-0.00688486791893184,-0.0116027359958535,-0.00135523267342008,0.000100218249234896,-0.00637047368061483,-0.00583667761465434,-0.0305998412437321,0.004944778001164
"1686",0.00224896683845155,0.00392181491631516,0.00519943025818548,0.00660320740980547,0.00387807076688973,0.00130691227267543,0.00218915198978031,0.00660488317782115,0.00117491973329531,-0.00302796768043412
"1687",0.00578755565574118,0.00597437559575842,0.0129308693731602,0.0111756233186944,-0.00666376801268831,0.00220999974396663,0.00982997269752572,0.00801940460271089,-0.0107182209356907,-0.0125284973465647
"1688",0.00446243123930445,0.00137028845312259,-0.0042552893374902,-0.00216226628832616,0.00826371061897957,0.00200320845864699,-0.000772625106166158,0.00699151233705009,0.000395436940975102,-0.0103806785639978
"1689",0.0115741924801478,0.0253194687163834,0.0307693876074153,0.0418974790548459,0.0123420725606518,0.012400427554957,0.0349463069816256,0.0277709823745171,0.0435572727272728,0.0217560449952168
"1690",-0.0016756824252091,-0.00489448259883574,-0.00497512576416059,-0.00531538450241187,-0.00590511261881532,-0.00345678635064461,-0.00388424535977672,0,-0.00196950996021172,-0.00380226857225308
"1691",-0.00699145163055248,-0.00558914930619414,-0.00833357676843305,-0.0223049373254478,0.00526941380453372,0.000991390717487661,-0.0172493392720627,-0.0112543001163529,-0.0287666110056927,-0.0091603372497493
"1692",-0.00462766383541002,-0.00382174228971155,0.00336147178951118,0.0035647438259363,0.00733906407825735,0.00376269805212459,-0.006410307420749,0.000236750347167414,-0.00320409505473651,-0.00731889206234926
"1693",-0.00235397863740894,0,0.000837388390326321,-0.00852462927033149,0.0107863069767165,0.00364976309253429,-0.00660496486358986,-0.00189658378360791,0.000862414719033699,-0.000388042802127453
"1694",-0.00289033913400416,0.00225677320406437,-0.00251048501437401,-0.00764280391353667,0.00205925886622804,0.00275194352160746,0.0034337169342562,-0.00237522603540463,0.00885155071748245,0.00155269384311052
"1695",0.0038454763866882,0.000675727816086491,0.0159397784293167,0.00409136733316218,-0.00700622373322946,-0.0021566258070751,0.00606639522000108,0.0050000521290976,-0.00776451630057939,0.00775195220958547
"1696",-0.00459668797803436,-0.000675271516339504,-0.00743171544691834,-0.0117447557139655,0.00244603548974598,0.00137533573511583,-0.00371050124234562,0.000236866172109274,0.00923389929388918,-0.00499997149863052
"1697",-0.00532827488197063,-0.00653007101696657,-0.00831980323791481,-0.0113996744022671,-0.0015016643620771,0.0016676837453109,-0.0100870138789952,-0.00213173278192802,-0.00612551751472812,-0.00425197135461264
"1698",0.0079162330004805,0.00770621140781746,-0.00419441397329035,0.0198725428457649,-0.00303366116302561,-0.00222613067040944,0.0152061794636764,0.00688366265922769,-0.0280074675928559,-0.00659936835062425
"1699",-0.000944564360772171,-0.0013493306453457,-0.0050545964920623,0.00384883927711432,0.00151192902091113,0.00167093866652879,0.000617431920802325,-0.00117870460813696,0.0198250427747024,0.00976938764059976
"1700",-0.00922119640445562,-0.0049550018956096,-0.00762078032119085,-0.00383408250975903,-0.00160444867719978,0.00137390308585239,-0.015431955732805,-0.00873274804405089,0.000944451455130668,-0.00154804612847681
"1701",0.00757684432811745,0,0.00170638162167713,0.0129898466627059,-0.000756476366934766,-0.00274385672606503,-0.00360491362177062,0.00309520362736482,-0.00511087435131308,0.00310081279751295
"1702",-0.00864507272610504,-0.00520598988512089,-0.0187392487930412,-0.00854881240631111,0.00406814493970686,0.000884172552361617,0.00440466934002237,-0.0113930750967044,0.00877262316266991,0.0069552021763386
"1703",-0.01164631663993,-0.0102389978888183,-0.00347218272720995,-0.0095808950953209,0.000282473234238356,-0.000490253794776851,-0.0114332352771741,-0.00384177943755915,-0.00188026482200143,0.00345352149477884
"1704",0.000725181168731437,-0.002758611459723,0.0235189501866695,0.00749685174929082,-0.00800573556914697,-0.00176899827654331,-0.000316891730980928,0.00964100462357553,-0.0101255963873533,-0.00726575415014186
"1705",0.0215576239688906,0.0205163592421747,0.0144679885132424,0.0235240200433435,0.00161385810468806,-0.00216461821729586,0.0239302807726354,0.0181426356770873,-0.0145904685227938,0.0127119685621264
"1706",0.00644300738833037,0.00609890410299641,0.0016780098753082,0.00445577105874606,-0.000284032740759499,0.00147881150440843,0.00959647218303439,0.00281367658351939,-0.0134384730048719,-0.00532534128258155
"1707",0.00399431561606867,0.0029186830341088,0.00167529267380817,0.00583720198870585,-0.00806007185874058,-0.00334789293786719,-0.000306800658162243,0.00327347949228995,0.00187605223288823,-0.000382403970200285
"1708",-0.00725410282023775,-0.0026863578995141,-0.00836135351936962,-0.00974938762015387,-0.000669405918622301,0.000197936220131867,-0.00322060976354099,-0.00838954737370112,0.00732720821741917,-0.00344303107689314
"1709",0.0139662277835269,0.00718296270725682,0.00927470317361445,0.00796990498618677,0.0125312955809564,0.00483993859709719,0.0181537473483555,0.00846052736886871,-0.00153561784040357,0.00767759687630321
"1710",0.00668296944943947,0.0147094110514143,0.00835425397668432,0.00627908016691703,0.00906932138561833,0.00570242945748234,0.0154126405424386,0.0139826347196401,0.0314068072575133,-0.00533326056285455
"1711",0.00675452697516055,0.00636924743820999,0.000828531702501412,0.000924406449227311,0.00215300490603765,0.0000973599548070858,-0.00193447581080408,0.00873360010287061,-0.00447339514163236,0.005744925346165
"1712",0.0000569647738586365,0.00152776093908602,0.000827845806006033,-0.00161596683082699,-0.00317603107926911,-0.000683768276922958,-0.00521833459326737,-0.00273424850036352,0.00102487191209888,-0.00228489091290041
"1713",0.00579177374428719,0.0126388582131125,0.00496280415398487,0.00971279598505248,0.0111528912734542,0.00694413171998853,0.0106414792783567,0.00525516453619557,0.0185855484662416,-0.00114502251469084
"1714",-0.00478891236411039,-0.00602535496065859,-0.0205763077918595,-0.0233620593927313,0.00389250504657435,0.00174839440073682,0.00207618579370772,-0.0065911371766455,-0.00502546791481284,-0.0152846645628761
"1715",0.00332228687738034,0.00736085799437491,0.0100843447829908,-0.00211087152869127,-0.00387741220001814,-0.00203609279998984,-0.000739910494803708,0.00205886833483948,0.00940237766100904,0.000388042802127453
"1716",0.00456763904170554,-0.000859718885829253,-0.0149751846146987,0.00470043600179837,0.00370746536743516,0.00174873702850697,0.00977478272244015,-0.000228267628651024,0.00431110874416207,0.00310321811263736
"1717",0.00159140306507433,-0.00408685625818384,0.00337824559949795,0.00584790574148597,-0.00341707121076229,-0.00096928575352373,-0.00689373326122233,-0.00411021443991255,0.000766449445307904,0.00386688312838346
"1718",0.00533383496388118,0.000647932793773176,0.00757578489335575,0.00325577895037621,0.00129725204543485,0.00135862990760027,-0.00841806008942092,0.00114627739346673,-0.00605081197994506,-0.00269645895743109
"1719",-0.00496701619415985,-0.00366934733842961,0,-0.00556323436797268,-0.00601499099759129,-0.00261767161576976,-0.00729820279735816,-0.00847423350418852,-0.0013099945654621,0.00308999375752017
"1720",-0.00283606601867847,-0.00498247146164232,-0.00501246350051698,-0.0102566356277185,0.00214141155942826,-0.00116661750194746,-0.00720181385320373,-0.00323415724267617,-0.0143519129158065,-0.00847131645656707
"1721",0.00238923122429258,-0.00631388509095021,-0.0109151624941681,0.00047117255416973,-0.0108240015177355,-0.00554654968388468,0.00634718120851163,-0.00324485058598456,-0.00618444506316651,-0.0124271349969011
"1722",0.00351847371011726,0.00591574834686903,0.000848738289412898,0.00612084047869321,0.000941407498666447,0.00196036855717185,0.00135179143579367,0.00279005913253672,-0.00110278852546963,-0.00432562145749138
"1723",-0.00316686893772888,-0.00936630081255219,-0.00848153907398208,-0.0201218915364818,-0.0119483121795858,-0.00449967282340402,-0.0151469905051396,-0.00765108198120901,-0.00197145338650662,-0.00276465649222335
"1724",0.00510569211051637,0.00945485785536548,0.0136868041614309,0.00310415356564997,0.000475953483275449,0.00304600141085198,-0.000152085276171943,0,0.00505688219116451,0.000792149946476695
"1725",-0.0126432713771688,-0.0154651244477736,-0.0185654870603837,-0.0180907312719836,0.00847058175136395,0.00264542270254764,-0.0121844265719044,-0.0135515048996323,-0.0081760457903155,-0.00712309554301804
"1726",0.0134913806996362,0.00553113969602781,0.00773880343691102,-0.00218200125104007,-0.0240656629186553,-0.0112371723940646,-0.0134132122217653,0.00450051367792437,-0.0149017512713459,0.00557991813609582
"1727",0.000169093359377648,0.00308012670014812,-0.00170662052036008,-0.00510204256035773,-0.00377157225607316,-0.000494224924520004,-0.000781468328420187,-0.000235952203057388,-0.00329897009413405,0.00435987023310913
"1728",-0.00203047986471128,-0.00592245222965404,0.0128205422736931,-0.00537252310939962,0.00465985811590719,-0.000889825624854623,-0.0034407590906389,-0.00165076852735579,-0.0114636793865259,-0.00670879114630474
"1729",0.0080244828987639,0.00441328218418136,0.00759493975953718,0.00171890438153932,0.00367113889195236,0.00415639123495937,0.00706232337070301,0.0011810070621312,0.00326664769130214,0.00437042702655299
"1730",0.0049896089004493,0.00241665063501451,0.00837517363615259,0.0161762766544939,0.00616088424659966,0.00482917927223059,0.00794755107784373,0.00802249942240563,0.0115588036069809,0.0043511245202319
"1731",0.00435085240917199,0.00416369333072764,0.0141195997064669,0.0190544826714996,0.00200918275260498,-0.000784543730002363,0.00247364737854561,0.012406456879863,0.000402373873075623,-0.00157540193747197
"1732",-0.00349919698429813,0.00240082820204801,-0.0016379717768038,0.00899410900166009,0.00601540525679334,0.00353345982661657,-0.00694019322760053,-0.00346825356780556,-0.0114221203346203,-0.00670606351599057
"1733",-0.0021737044679947,-0.00239507803116468,-0.00574235289307712,-0.00609900021755327,-0.0075929311418903,-0.00371674294022262,-0.00760983767451107,-0.00719252347705712,0.000406794134958588,-0.00158862234773016
"1734",-0.00312776074299592,-0.0104758462156667,0,-0.0136887912903608,-0.0170236353211621,-0.0054981847205644,-0.00876370254352765,-0.0100492354256175,-0.0230174385445491,0.000795534102772777
"1735",0.00806840983439305,0.00992518059062131,0.00412538316889766,-0.000957256541302076,0.00165366062350758,0.000888848922883323,0.00536783166580457,-0.00165205656538103,-0.00149850978608446,0.012718632235597
"1736",0.0050027838754414,0.00502294451394891,-0.000821631645000265,0.00718547473846298,0.00932551065031872,0.00286051876249083,-0.00298349683016108,0.00118192037635145,-0.000166783388914737,0.00313971495238485
"1737",-0.000995599065921282,-0.00173881151358657,-0.00740143324569009,-0.0128417656959399,0.00288681034124316,0.000786782644772277,-0.00425270689540158,-0.00661307673897971,0.00450301041532697,-0.00117365263192004
"1738",0.000276745141073675,0.00152401037830718,-0.00414228735851108,0.00337275796882852,0.00374261864468628,0.00216142927350926,-0.00284722585389663,-0.00071316691543144,-0.00531295870258142,-0.000391771302957644
"1739",0.00243521407461333,0.00369497399535801,0.00415951727433406,0.00648237800359341,-0.00172117735032051,-0.00225487374739031,0.0103108633505191,0.00499634605324895,-0.00300451510599231,0
"1740",-0.000662560746611085,0.00346464723404005,-0.000828346125503643,0.010257640480057,0.000287395489634079,-0.000589495805829343,-0.00926369217225087,0.000473633823036002,0.0103800268741003,-0.000391844188296631
"1741",-0.00259663178722014,-0.0079842991874709,-0.00248756288208019,-0.0210152000158139,-0.00777804520347336,-0.00429479459109017,-0.00522982459092292,-0.0134881818142905,-0.0258491721420673,-0.00117599337105756
"1742",-0.00432039075458268,-0.0100067652899865,-0.00415633920220759,-0.00337671226310399,0.00367730647208875,0.00178076214796707,-0.00111517075820333,-0.00407763962492658,0.00323181658051008,0.00588701097795474
"1743",-0.000111609234185295,-0.00549335608859336,-0.00751238321490977,-0.00121016006670971,-0.00954554543235175,-0.00454211386074455,0.00223289375963254,-0.00192673157224277,0.0169549001098246,0.00195089246041613
"1744",-0.00439567634369042,-0.00397690059229394,-0.00841074462559011,-0.00581531204420715,-0.00282341759058113,-0.0024803750301523,0.00111392846847846,-0.00506748159894321,-0.0138379127529001,-0.00116836855358804
"1745",0.0111772372072401,0.0135314221356588,0.0127227716976346,0.0221788830733984,0.00478392266199323,0.000895158961147891,0.00778909195794864,0.00654847818282422,0.00211327129044969,0.00350880445250534
"1746",0.00254220159083851,-0.000437775712838429,0,0.00143073554758044,0.00233186216319448,0.00119219831136164,0.0064668196672637,-0.000963985748440144,0.00986923635927694,-0.00349653579214948
"1747",-0.00358317196666069,-0.00394098392704456,0.00167529267380817,0.000476137435551971,0.00717360912137921,0.00416778192522482,0,-0.00241175304635033,0.0175409203346064,0.00311894620786823
"1748",-0.0112308702458949,-0.00681473620294459,-0.00919757549004374,-0.0221324767682349,-0.00769978184181841,-0.00385424431188808,-0.021626763034379,-0.015957641970949,-0.0078804711869972,0
"1749",-0.00330141558947161,-0.0108456533845702,0.00337572568024869,-0.0058407870831042,-0.00378266840566888,-0.00287685366390855,-0.00672733876404819,-0.00491350586573314,-0.0212642725362876,-0.00932762588406888
"1750",-0.000112035621518625,-0.000447653606258203,-0.00841074462559011,0.00244808127722829,0.00486778321443193,0.00149278345021919,0.00403147452006758,0.00197486599288199,0.0092146080884723,-0.00392313431467806
"1751",0.0062316550954935,0.0123125512826749,-0.00593700848248901,0.00659341703933958,-0.00368158208041103,-0.000497317339381742,0.00112405465680498,0.000246557438666972,0.00259679182267036,0.00315080387494393
"1752",-0.0031803633823827,-0.0045769927623448,0.000853202755772831,-0.00873393212545215,0.00447345004770572,0.00318084602745894,0.00529457852568549,-0.00813011005727615,-0.00868911339812661,-0.00471136123717364
"1753",0.017072588380773,0.0156249711304819,0.0195842586644444,0.019904401460036,-0.00503473207815341,-0.00376545445357379,0.0175552092808595,0.0116743143901157,-0.00876528430231294,0.00197235968110299
"1754",-0.0011557120434833,0.00307708334971979,-0.00842457093754201,-0.0184021120824279,-0.000972679076311822,-0.00417682369817651,-0.0122334368567517,-0.000491192947463137,-0.0237224808798361,0.0023622536040393
"1755",0.00581711283321074,0.00328648133101139,0.00339848254329822,-0.0014797844103045,0.0153891285733074,0.00309615444678157,0.00778020637570975,0.00326201663633063,0.00975441560703727,0.00785547348507354
"1756",0.00534231714254618,0.0109193715140758,0.00931409646758241,0.00741100657865013,-0.00565961436017193,-0.00318656993131339,0.00141526883978504,0.00825438623348229,-0.0031913230431031,0
"1757",0.00219162432380093,0.00691293203622867,-0.0134228427306087,0.00588529835676277,-0.00800687155879154,-0.00389483392492573,0.00174712828339629,-0.0017367025842262,0.00458594791035738,0.00311765026524369
"1758",0.00508367787780228,0.00493433728424875,0.0161564666841152,-0.00853255643227091,-0.00385363015966578,-0.000863428782049702,0.00110950756268147,0.00372793502720858,0.00551248932838044,0.00155406033549488
"1759",-0.0000544121886295601,0.00533758475219037,0.00502097315992245,0.0154906118006393,-0.00284076354957374,-0.000603869420534586,0.00126667915505285,0,0.00325513968228774,0.00271524598323292
"1760",-0.000162846482962831,0.00339761564084018,0.00915889833425232,0.00435819431998996,0.0068756769385343,0.00271627128134089,0.000791065387079959,0.00940803070394436,-0.0147712086380325,-0.00580270831542484
"1761",0.00473274427585668,0.0042328447711486,0.00165018245851822,0.00771492186332634,-0.00634037427075351,-0.00451423844713095,-0.0031605177829771,0.0105468354667746,0.00632640615587476,-0.00155639897877735
"1762",-0.00958357233229357,-0.0229714769032681,-0.0164743637417133,-0.0385169086798963,0.00304287219462873,0.00393017080662283,-0.00158552460259553,-0.0189319443849404,0.0161901218690117,-0.0144193330254777
"1763",-0.000163962600562395,0.000862910208264012,0.00586266128282431,-0.00174171934489242,0,-0.000602423194756896,0.00587504900718172,0.0054427189813,0.0109322118644068,-0.00632664688813733
"1764",-0.0028981502826646,0.00172420130060025,-0.00333059262377777,-0.00947160256978363,0.00420912203177903,0.00281214899598115,0.00410410682125573,-0.00344440640572108,0.00176040739575489,0.00119377599891823
"1765",0.00614197965793539,0.00709968572422426,0.00417719960614549,0.00427764127835983,0.00253377639152919,0.00160250441633503,0.00345851167049349,0.00172841592467576,-0.0056903765690377,-0.000794901731337117
"1766",0.000217787133558911,-0.00170920349666004,0.00166398013923241,-0.003257170043795,-0.00272210793774041,-0.00489988753076087,-0.00156655176210463,-0.00419074961796062,-0.00589123884867859,-0.00954649111203931
"1767",0.000653799927067933,0.00085615610940093,-0.00332245489836314,-0.00527909980758179,0.00584872173028916,0.00261281111526857,-0.000470919335393338,0.00173276452052984,0.00287839477958696,-0.00803205995609246
"1768",0.00272289510526758,0.00962157149254539,0.00666680607419434,0.0176902124957989,0.0119211967084203,0.00841853121715275,0.0119310914806998,0.0071658313116485,0.015195027985776,0.00647764372042814
"1769",-0.0133050490784556,-0.00847106664120068,-0.00662265412345686,-0.0119195213805291,0.00498075997391956,0.00288210416723511,-0.00651574782207143,-0.00662411011825814,0.00631959909663071,-0.000402247119002164
"1770",0.0108976041658873,0.0128149500271262,-0.00249997991095841,0.0108068352985771,-0.00457472739924614,-0.00376578548176321,0.00624618218694972,0.00419868390632216,-0.00933728332516814,0
"1771",0.0053900633065993,0.00421767010813356,0.00751873642288836,-0.000248631436483904,-0.00105302979862298,-0.00089507510028386,0.00465544716043365,0.000245436390118314,-0.00191838353422624,0.00281690432515114
"1772",-0.00129961423311564,-0.000209866158304872,-0.00331660017421287,-0.0054713097231931,0.0067087852402461,0.00278840221301846,0.00231702680191215,-0.0012292651351844,0.00108638639189751,-0.00160515579427789
"1773",-0.00422965280296661,-0.00483097740867555,0.00249588929282929,-0.00500131582988528,0.00418847114298515,0.00238216633380683,-0.00323633486581232,0.00221580881069516,0.00951664571736677,0.00120581268813291
"1774",0.00294049879368719,0.00548744788815414,0.00165967593978622,-0.00150791013280804,0.000758628944358186,-0.00108977098140151,0.00695726960445597,0.00343903584791239,-0.0101711982138428,0.00240863827526017
"1775",0.000651737163044119,0.00125933269624867,0.00248541199249908,0.0133400175901908,-0.00246315387371476,-0.00277611838178082,0.00261034382461078,0.00416164771635552,-0.00426060996476041,0.00480578379051
"1776",-0.00819324062110605,-0.00167700686925909,-0.0198347351902687,-0.0245902616386336,0.0141499949736412,0.00676171991182906,-0.000459498359341892,-0.0107266606576381,0.0218139018069652,-0.00079720148395801
"1777",-0.0213361875474329,-0.0317094472823241,-0.0151769208364022,-0.0262284166879168,0.0064613882291602,0.00404914242410381,-0.0147080211098678,-0.019713935913466,0.00410542734128061,0.000398959814302602
"1778",-0.00491899036481624,-0.00542187618632173,-0.012842622763293,-0.00392278956382464,-0.00697764688974145,-0.00304967103621756,-0.00606437293748829,-0.00351936432901567,-0.01087580332917,-0.00677829885603132
"1779",0.00595460367741385,0.0109029725372831,0.00867309413191708,0.00630090085560919,0.00243599612781376,0.00147987569817087,0.010168640630309,0.00983867282343742,-0.0000826884927470628,0.00481735918529047
"1780",-0.0096048501926338,-0.013805092939951,-0.000859806438417321,-0.0143490432485732,0.00822501541619491,0.00472918334842221,-0.00464607531538297,-0.0102426433947256,0.0125672099024525,-0.000799030209567286
"1781",0.0106002524797748,0.00393705347119444,0.00172099702462947,0.00926430586431071,-0.00287425991687129,-0.000980235939280205,0.0121364181033763,0.0070672969896397,-0.0220462478807361,-0.00399842815131779
"1782",-0.0058583624171209,-0.013725635276889,-0.0266322266006417,0.00157343527344356,0.00669400989847424,0.00392605391050815,0.00307438232051815,-0.0105264103327246,0.00267177931047291,-0.00120436045501515
"1783",-0.0225053570790749,-0.0203224151897203,-0.0203000320639,-0.0282796243160389,0.0121846658340359,0.00543587796797351,-0.0145591698737543,-0.0167173142460026,0.0102423519108119,0
"1784",0.00700491829914873,0.00901914214811605,0.000900685013299318,0.0202102238519306,-0.0106109403483193,-0.00301952476164769,0.0104200244061698,0.0118495333213144,-0.00272009561490272,0.00763659306640951
"1785",-0.00125463522405989,0.00402236586881988,0.00180027428201068,-0.00369778731856263,-0.00924566259974591,-0.00361561248378184,-0.000308265142624942,-0.00152750368888532,0.00247956860037313,0.00199447064194791
"1786",0.0131873955763431,0.0213665740493796,0.011680392242144,0.0209436117180177,-0.00429242642467176,-0.00186279709457948,0.00739062213461383,0.0137684572353425,-0.00041225986963267,0.00398087837775551
"1787",0.0123953789777134,0.0124211904714726,0.015985560842982,0.00571274756391049,0.000843315305525838,0.0026522275638341,0.00672456029474455,0.0125755490288733,0.00767073585732003,0.0114988169728101
"1788",0.0018368770817585,-0.00258302744482708,-0.0043707241351677,-0.0111023982141404,0.00280934546416844,0.000490120937892913,0.00910907504345926,-0.00571264288894069,0.00613898675843472,-0.00548796906493509
"1789",0.0109439382033836,0.015106002467858,0.0140475597788472,0.0216710469282888,-0.00578983653422227,-0.00440716865563273,0.00346011427117521,0.0174868516757807,0.0117149611408225,0.00512409213369813
"1790",0.000494422287936613,0.00276342536185781,-0.00173161993776583,0.000255646380447727,-0.00516562633528284,-0.0023606316752981,0.000599805026646694,-0.00147367580602142,0.00056287390991594,0.00196075756439518
"1791",0.00516292145019803,0.0067840680026392,-0.00867292542234221,0.00102196791643006,0.00566498668593929,0.00473284957760645,0.00389564232921757,-0.000491408879728317,0.00851882986418051,0.00547949829681849
"1792",0.00551862479270682,0.00547445489345177,-0.00437435294530097,0.0122511540860588,0.000563270978675368,-0.00068732013761208,0.00402970882141251,0.00369005794983024,0.0132281777548517,0.00350334094595328
"1793",0.00119551665435313,0.00607365460065346,0.0219682261848091,-0.00932955102590438,0.00225123975639185,0.00245522464499559,0.00594628857915591,0.00955870563112704,0.00196618164425977,0.0143521342519306
"1794",-0.00662157851679224,-0.00666120869494935,-0.0120377441263446,-0.00687191957534572,-0.00421243838949537,-0.00195900823757589,-0.00029539409233148,-0.00242756035370528,-0.00886974083406999,0.00267682779140133
"1795",0.00590101290795109,0.00586756030076185,-0.00609246245569717,0.00358809702688911,-0.00244410252247829,-0.00108030244853619,-0.00177403153725875,0.00803129860201968,0.0105329930434701,0.00190703312623652
"1796",-0.00114084861125441,0.00166675348202716,0.00788094543605022,0.0068945229440196,0.00527751730538784,0.0012779728570218,0.00162884701793442,-0.00193173865198537,-0.000156708466406141,-0.00266463921158044
"1797",0.00554680657468443,0.00665546443155329,0.0112944766599865,0,-0.00253083464561277,-0.000981535322705285,0.00162650311036061,0.00241912589262228,0.0110519123522197,0.00419845517025497
"1798",-0.000378679076319499,-0.000826439047680649,-0.00343617605926005,-0.011412553422717,0.00892811103873514,0.00343819058106498,0.000442653484744593,-0.00241328784550887,0.00170557400939697,-0.00456098027062002
"1799",0.0000543035174882522,-0.00475605571554316,-0.00431050921478993,0.000769741452186778,0.00530998862149223,0.00293679880250863,0.00280314452440567,-0.00362850186583852,-0.00851331894131058,-0.00267273931650935
"1800",0.005247519420994,0.00540214090144975,0,0.0189692045648193,0.00546688743966817,0.00117138622202329,-0.00102978076511995,0.00194221887750778,0.000702490042131743,-0.00306282394495516
"1801",0.0025291764572426,0.00289303364913129,0.00519476357476401,-0.0067923961971631,0.00055336520674576,-0.000974702766191271,0.00662710918396803,0.00508847148213265,-0.00452413427123555,0.00345609488391885
"1802",-0.00703197854851101,-0.0247271095696143,-0.02325572433529,-0.0177304239175949,0.00667511246483787,0.00494553679680654,0.000731675867590598,-0.0106073005763221,0.0209214068111252,0.013777356550581
"1803",0.0140556868394459,0.0202833311219377,0.025573190273394,0.0170190410816353,-0.0150414998691766,-0.00768392018064179,0.0122808341707927,0.0160818578278172,-0.0123570503223529,-0.00377495795619198
"1804",0.000906192250986981,0.0012422807409278,-0.0111780332644545,0.000760852182728255,0.00214177199076415,0.00107808479297744,-0.00129984917877157,-0.00311750086318274,0.00163200195387003,-0.00833649397690217
"1805",0.00229024590615245,0.00868681222070644,0.0191305150499117,0.0141878706003222,-0.00984933277386657,-0.00430812847657558,-0.00477221131328798,0.00793842742354545,0.00993094118962645,0.00917079873772564
"1806",0.000425066937856489,-0.00676639601498608,-0.00682610462198219,-0.0127404490971441,-0.0062880011237002,-0.00432667947218113,-0.011333873391231,-0.00119354764487245,-0.00829685808245906,-0.00454367128187516
"1807",-0.000530972462193469,-0.00639971424700048,-0.00429543493654161,-0.00683192567828306,0.00141677085222103,0.00108585745481871,-0.00367413687991902,-0.00931915098388647,0.000309931065455959,-0.00836828159099012
"1808",-0.00494274612910206,-0.00498642623452172,-0.0103538379914746,-0.011209847248683,0.00264033191373736,0.000987215451853762,0.00545782539594675,-0.00651217015991012,0.00565318649217117,0.000383577422433889
"1809",0.000267231362070852,-0.00292362001099078,-0.00959009465783645,0.00206095561562214,0.00696021058173102,0.00394214857813036,0.00220082423251378,-0.00534090572942103,0.0146310949127437,-0.00268401243046767
"1810",-0.0112132832895925,-0.0215704969635806,-0.0167252577314165,-0.0179994392402063,0.0134500207576576,0.00589038240491258,-0.00322072173650334,-0.0126921934530783,0.0034153917507358,-0.00461366569400934
"1811",-0.0028081011204566,0.000856235097046021,-0.0116385617594372,0.00549864595983962,0.000184607549674087,0.0000976029493193753,0.00029357199440927,0.000741278331982009,0.00673170677617474,0.00540753876743816
"1812",0.00904371279496163,0.013045197417576,0.0108696552313836,0.0122397145220519,-0.00746401945443931,-0.00400105350395552,0.00161512785768059,0.00914059055659777,-0.0109692481907178,-0.0111410364454776
"1813",0.00713765280928746,0.00865529510360208,-0.000896216165984676,0.0138924329743357,0.00362040167464595,0.00244911410661386,0.0043975695695615,0.00538542700150724,-0.00774843518496227,0.00505051615747321
"1814",-0.00532857651758678,-0.0146503799461984,-0.00538082455566069,-0.0213142973445669,-0.0077702939349944,-0.00928548914995786,-0.0176592307987379,-0.011200226609252,-0.019369155541615,-0.000386463282109228
"1815",0.00583943694332167,0.00127431191590754,-0.014427435739676,0.00440755166262297,-0.0017714010617651,0.000198085760654498,0.00133719697667534,-0.0123125040597395,-0.00179557348100801,-0.00464046671164819
"1816",-0.0038787425882586,-0.00318190603716972,-0.00457476529907697,0.00619506057432218,0.0108340101822562,0.00187360614903342,0.00816017300369265,0.00170640105365072,0.0047708430723381,0.000777070152832904
"1817",-0.00413518315486194,0.000212861183034097,0.00367650936961517,0.0097487269024279,0.00711455834726893,0.000394000369787983,-0.00588642146259388,0.00325668833618198,-0.0178251808373535,-0.000388273345873769
"1818",0.00474568005392295,0.0129787645127637,0.00457892993943276,0.0114330543442056,-0.00376139132089237,-0.000590516494081039,0.0073222108040647,0.0099875607420099,0.0018228245363765,0.00660197167429399
"1819",-0.00719199951459715,-0.00189047028350231,0.0072924889441075,0.00226084516403802,0.00782769387818494,0.00423434545557688,-0.0111490997127036,-0.00494455323488718,-0.00791076630295806,-0.000771634106060737
"1820",-0.00210849801743918,0.00273569195528633,0.014479588304168,0.0130322306445811,0.00502492545898914,0.000980445332549928,0.00481056091134091,0.00993793443923807,-0.0065386171265891,0.00888022757835838
"1821",0.00492997473861312,0.00629600593100221,0.0107047164887593,0.0079171268547078,-0.00563666178690281,-0.00352650843013691,0.00658298272882218,0.00984000633684512,-0.000240773745590395,0.000382775466384988
"1822",0.00819417148655854,0.0068820319668268,0,0.00662710685299617,-0.00246845934348705,0.0000984803402415135,0.00579663258132546,0.00292342431103254,-0.00762682253736069,-0.000765021771425012
"1823",0.0066310466328583,0.00683537151654967,0.00264791451346813,0.0117044699123805,-0.00854602871834431,-0.00206827394584141,0.00635440643421736,0.00218604992530369,-0.00177980744454487,-0.0122512563764504
"1824",0.00334654099378606,0.000411133797732388,0.00880298223549691,0.0019283634068965,-0.00574657799987055,-0.00434204580403341,0.00014676850026496,0.00799799845295013,0.00753708572442724,-0.00232554975998711
"1825",-0.00132335242619919,-0.0026731487871432,-0.00523582566358893,-0.00384899648218173,0.0043814873786856,0.000693319917830948,-0.00352357362813194,-0.00384710978440939,-0.00321751930501923,0.00815851687320612
"1826",-0.01182262223015,-0.00371138308572283,-0.00438596223945109,-0.00265643589916253,0.00668254777725119,0.00614152363218823,0.00397818745256528,-0.000724076720451383,0.0133150583168988,0.00462429368806183
"1827",-0.0110512924602513,-0.00393211022232531,-0.00969165830082752,0.00435819431998996,0.00599291907438881,0.00236258772069253,0.00102713168725943,0.00458936697043333,-0.00525600063709475,-0.00230146453460378
"1828",0.0041228871968797,0.00332437689146459,-0.0213521424803965,0.0115719626014283,0.00238284197941385,0.00137516511498759,0.00557121741997557,0.00264467814297542,0.00944673734859536,0.0115339861699637
"1829",0.0107507728593821,0.0132533472788476,0.0145453020511472,0.00762644482578789,-0.00493685233297969,-0.000294539402566296,-0.000729027278845273,0.0115111211565668,0.00182412568242118,0.00266054900521828
"1830",-0.0210057543878807,-0.0183937347545238,-0.0286738127239887,-0.0106434488604318,0.00928043686911839,0.00421890423019944,-0.00889988530797681,-0.0113801231798667,0.0054623337555415,0.000379147925316126
"1831",-0.00900889097911906,-0.00666249520458839,-0.00369007559010015,0,0.00810265586281189,0.00205128425318191,-0.00603553159610304,-0.00167836125132892,-0.000629887400521389,-0.00454719271475734
"1832",0.00787859654570622,0.00482095433377272,0.0138889835912086,-0.0021514456631494,-0.0026191693640516,-0.00155966495364668,0.00370241048129238,0.00384354705405276,0.00724807374143221,0.00913592825592224
"1833",0.00688764320268742,-0.00438063979792325,-0.000913302290496132,-0.0150935091978086,0.00624791233344291,0.00117163128546882,0.0106239792952638,0,-0.0184591320838347,0.000754344303005805
"1834",0.0104776667967832,0.0111042090548261,0.0191954327890091,0.012649106117266,0.00125968925594022,-0.00156068201577608,0.00598651947878159,0.00885363653552962,0.000398462035197555,0.0018846720080643
"1835",0.00139687062334226,0.00580180482041293,0.00269066150546138,0.00912774146044026,-0.0109642413281056,-0.0056655562766359,-0.00275772114478223,0.00450656969896723,-0.00629282295449407,0.00225738301863121
"1836",0.0034871736240023,0.00185407462446618,0,-0.00618875600715763,-0.000817976808664578,-0.000196624514936183,0.00422063300518261,-0.0028336848087227,-0.00408819238476954,-0.00337844807662935
"1837",0.00454444647817831,0.00658049371349945,-0.00715551198374254,-0.00263457994089977,0.00336506712685103,-0.000393092628904967,0.00333314131494133,0.00497291645215991,-0.00370250327917743,-0.000376565178978328
"1838",-0.00234177648601708,-0.00326878668920683,0.00270258077537555,-0.00720496925608372,0.00570969907986307,0.00255576726370244,-0.00303317527169888,-0.00282734659238848,-0.000161552756192895,-0.000753569186683123
"1839",0.00202729099560206,0.00143475767135781,-0.00359362882157621,0.00096766619864419,0.00189259362642935,-0.000293775383746531,0.00333230471087487,0.00307173414320649,0.00646409168610051,0.00603313866066468
"1840",-0.00819860115448257,-0.00450259648759155,-0.00631210806478155,-0.0135333035042509,0.00143918025083822,0.00137286557531402,-0.00346571577001165,-0.00494701129744535,0.00698460191047867,-0.00412292080413723
"1841",0.00316706395104394,0.00328921955294637,0.00544450120457962,0.00489985249858726,-0.00485001168702304,-0.00146916912685713,0.00521683775742043,0.00378784297637869,-0.00438493980706378,-0.00338731004097692
"1842",0.00465519969835326,0.00840176722398067,0.00270748448299618,0.0095075730064198,-0.00135387792932329,0.000882694015244434,0.000576528134822896,0.00589618323064234,-0.000160121720694795,0.00264346846756669
"1843",0.0029827437254204,0.00792524878257073,-0.00270017380431964,-0.00193189215884337,0.00415774467637142,0.00264565785333182,0.00446621164268324,0.00140699096014196,-0.00512574078867745,-0.00527299793137248
"1844",0.000105961544206501,0.00201618514201152,0.0126354124714783,0.00120965728569833,0.0107278198490377,0.00287983983463014,0.0077452558489215,0,-0.00338108192415798,-0.00757290238187724
"1845",-0.00143362224723276,-0.00321926325385102,-0.00178245093244578,0.00555818920358297,0.00615939783755781,0.00146454947379171,-0.000426841795685529,-0.000234016452356878,0.010177665343029,0.00267073913185523
"1846",0.00191433366264304,-0.000202002738843632,-0.00267845060544758,-0.00552746649896529,-0.00603295636562529,-0.000585194580422499,0.00355967102906374,-0.00117127176248477,0.0092755718739097,-0.00228319130765142
"1847",-0.00870389321444054,-0.00222078329441677,-0.00268611665464968,0.00459176736415667,0.00401708458694916,0.0011707435618038,-0.00368912829374934,0.00422054727351795,-0.00190142606638066,0.000762844652970829
"1848",0.00588936979793631,0.00364219362181983,-0.00448795430549931,0.00529233871672186,-0.00355646915908048,0.00077985844817241,0.0116777874875449,0.00817183361863894,-0.0143673992451008,0.00266768573702603
"1849",-0.00106460960087595,0.000806616399431359,-0.00360699048728552,-0.00239310095578893,-0.00428265043456733,0.00107095924307798,0.000563262178318036,0.00115779908357183,0,-0.00304070567216974
"1850",0.00149202242802016,-0.00423054446729654,0.00814455466051633,-0.00167916405356994,-0.00322590515145038,-0.000778505065291979,-0.000140884185418466,0.00277577564208276,-0.000563743264294869,-0.00495612882897922
"1851",0.00973608485200028,0.00809222997721504,0.000897700619699515,0.0168190184012256,-0.00404520258288432,-0.00262845202718753,0.00211047636753481,0.00553631292060053,0.00676876723237352,0.00229889807629657
"1852",0.000895829029729178,-0.00220760835596256,0.0134531081452025,0.00378067447814767,0.00866551850326314,0.00390456637774994,-0.00589711404346149,0.00206500692409173,-0.00272133819879405,0.00458713250180853
"1853",-0.00473800636800326,-0.00140789646640893,-0.00530979013890354,0.00706228068507841,0.0108271328075202,0.00456906609868635,0.00254239898087327,0.00251826289632739,0.00971107559728845,0.00456614763446561
"1854",-0.00878024116566489,-0.00382677900443196,-0.00978653049391653,-0.00935047533273758,0.00796738167568178,0.00358119100332743,-0.00169071218753047,-0.00159867070798481,-0.00826644159075485,-0.0060605625859117
"1855",0.00346837323111826,0.00141529746411817,0.00179686434587989,0.0132140821747351,-0.00281054858701446,-0.00212183028855228,0.00733847363036033,0.0036596817870469,-0.00216395773416589,0.00114331630053921
"1856",0.00366934160693488,-0.0014132972281351,0.00179404017978091,0,-0.00739813048070015,-0.00125618480499179,-0.00364220287019634,-0.000227967682430719,0.000642586345381391,-0.000761353473580639
"1857",-0.00630486114184736,-0.00545893418645294,-0.0116385617594372,-0.00815103465420963,0.0022183250518637,0.00290269906423712,-0.00309356946991968,-0.0093459098081653,0.000882966754166548,0.00190477512353748
"1858",0.00842435789636764,0.00833505423851855,0.0117756129581053,0.00774820996777037,-0.00610876606602995,-0.00154380292090195,-0.00394923661081603,0.0043720889287,-0.0024059908187346,0.00190111471928089
"1859",0.00243210569196428,-0.00100810484192193,0.00984756024898625,0.00698998976828369,-0.00142557409959776,-0.00106253308740156,-0.000849602294238361,0.000916291622828469,0.0022509767847172,0.000759081054928057
"1860",0.0040086228791576,-0.000403629203857725,0.00975170390417501,-0.00185095981354844,0.00535249761452072,0.00203128405798969,0.00751121685079537,0.00595095456184991,-0.0012833560805865,0.00227528168495428
"1861",0.00614680432246706,0.00868153200279176,0.00790180117082673,-0.00857695793699642,0.00585626380366211,0.000289431475011037,0.00604876202989724,0.00227531542174408,-0.0213637776666328,-0.00832387743504726
"1862",-0.000731008768030117,-0.00460347290802909,-0.0043553013201435,0.0058453568458916,0.0123500043767188,0.00550077102293622,-0.00405514336404755,-0.00567520094380325,-0.0053344358692563,0.000381450015833007
"1863",0.00517275376438819,0.00361939135087241,0.0113737212407337,0.0027894961139745,-0.00531541961334747,-0.00124721229545122,0.00126369588313135,0.00525082459263859,-0.00214517332042496,0.000381422326485303
"1864",0.00161140961069961,0.00140273193959461,0.00173002545133616,-0.0136767991553192,-0.000438049842369503,-0.000769077123965789,0.00490729687626401,0.00272584925121921,-0.00421698355850864,-0.00762479245482162
"1865",0.00114173566134701,-0.00080038611816835,0.0120897433719218,0.00305540786984704,-0.00743364353466069,-0.0045760873633206,0.00181431994101477,0.00385042113605616,-0.00606163746574784,-0.00115257963929916
"1866",-0.000518271890949329,-0.00300379734154399,-0.00170650244485182,0.00562319162863911,-0.0123050687087572,-0.00503239057733507,-0.00125366316603681,-0.000676861277936425,0.00258984968896869,-0.000769141123897699
"1867",0.00202286835461418,-0.000803269484785929,0.00683758328943318,-0.00559174815721208,-0.000269165639715463,-0.000777875595455502,0.000976121533466268,-0.00293529386561886,-0.00208315970197215,-0.00269442259198116
"1868",0.00652202505082089,0.0082412323177059,0.00254673956756557,0.0105436987028025,0.000448339116790208,0.00145996941779258,0.015603371285063,0.0040759455279189,0.00751504663468516,0.00115791773421514
"1869",0.00478252371772392,0.00737640407351225,0,0.00996976117144732,0,-0.000777346255189326,-0.00205784679035392,0.00902117849876727,-0.00041441238473694,0.00424041755856797
"1870",0.00102401168073785,-0.0017812250448721,-0.000846701817121764,0.00367315893108522,-0.00143371556394933,-0.0014594692199198,-0.0107215975830461,-0.00447005935350731,0.000331655747187964,0.00422274939862954
"1871",0.000102372843471255,-0.000792821514258635,-0.00847464073402759,0.00526070086067754,-0.00367976605854115,-0.00175344565447144,-0.00514094158383271,-0.00202102427028594,0.00613341887884933,-0.00267588302880972
"1872",-0.00347679105334142,-0.00674611718950113,0.00256398685324943,-0.00341292822679806,0.00180191439947341,0.00136601648044854,-0.00405032783066739,-0.00517372854534892,0.000164799408228111,-0.00268298369309872
"1873",-0.00707967230354967,0.000199709911202106,0.00341019046823954,-0.00479457940259254,0.0089007852417915,0.00389825734554972,-0.00294484442777754,-0.0027140407520081,0.0101309196892869,0.0142198340612605
"1874",0.00304852073534434,-0.00139798198335928,0.00509757035047498,0.000458925501217955,-0.000534396883402954,-0.0019414339656878,0.00253133101969172,-0.00385513565577,0.00260926290451113,0
"1875",0.000823871442128477,0.000199876524511922,0,-0.00458637715612165,0.00249680727605073,0,-0.0050504869914515,-0.00455267149096272,-0.00439168025692638,0.00303140980953276
"1876",0.00277973586695057,0.000199909603764148,-0.0016904705148022,0.000230467794213762,-0.0079162963980921,-0.00418283101046546,0.00112835896312591,0.00114352494525938,-0.00114359583636003,0.00113334305133139
"1877",0.00733969111532917,0.00799675711313763,0.0135477937928126,0.0110548205255547,0.00771045654175029,0.00527439914251215,0.00619705908389512,0.00776599061653838,0.00318939322202638,0.00415104216286699
"1878",0.00112099603006,0.00238025321977342,0.0175438808281159,-0.00569452510407553,-0.0128118332795281,-0.00252596776919467,0.00769856156708637,0.0031732692284443,0.0348088698917237,0.00977074474588324
"1879",0.00203008700161322,-0.00257231789976309,0.000820889750491105,-0.00206203284584783,0.00757065081889774,0.00116896372772257,0.00347305299332867,0.00247021474684139,-0.00346622020692899,0.00186078579704874
"1880",-0.000306164558413702,-0.00178536871790413,-0.00820341823720949,-0.0020660001830991,-0.00313042696737253,-0.000681233852281915,-0.00235329191845324,-0.00547574519332217,0.00276678260869567,-0.0037147358734172
"1881",-0.00602431330255515,-0.00765390629373208,0,-0.000460192321684594,0.010138938918119,0.00408938728444075,0.000461848721070357,-0.00183517144763723,0.00102487191209888,0.00149140393515124
"1882",0.00451998480319959,-0.00123380621722002,0.00349792784384628,0.00211113081164682,0.00257578628877853,0.000969757058827403,0,0.00666501669400565,0.0000787131813189124,0.00148918296182177
"1883",-0.000715782115099706,-0.00144147504885517,-0.00331956001170719,0.0011571520327136,0.00478443897340419,0.00261548372224052,-0.00111906712686571,0.00616444477671907,-0.00204736596657007,-0.00408908711055656
"1884",0.00194435332542864,0.00123721141439415,-0.00249796214402431,0.00231197568217945,-0.00149890474757186,0,0.0060206540266603,0.00476504732637251,-0.000552347497379868,-0.00186641921430597
"1885",-0.000510851744507379,0.00041198371673179,0.005008435169503,-0.00276781177135377,0.00247245390214057,0.000772929670739053,-0.000834913107829793,-0.000902991409806653,0.0108952230887345,-0.00598361722093199
"1886",0.00669342625291303,0.008853099318052,0.0174415461942337,0.00948400392210913,-0.00837243819230082,-0.00326924796312866,0.00250711395741776,0.00565069902597792,-0.00265538908612728,-0.00300977948909364
"1887",0.00101489873954819,0.00102050054741532,-0.00244875275584389,0.00595768063068935,-0.0106876737614684,-0.00407592582032568,-0.00111137308991638,0,0,-0.00188676673158761
"1888",0.00491816024214886,0.00550433594371369,-0.00327337986748066,0.00592258070818752,-0.00360086286252326,-0.00204593575228884,-0.00472961919936621,-0.00134858969476326,-0.0042286062074065,-0.00189041117318534
"1889",-0.00348152429795245,-0.0115570001875882,-0.00738920202197157,-0.000679078072414518,0.00731819774121178,0.00244153577684458,0.000978632193323614,-0.00472615854899971,-0.00110103016354102,-0.00795447621105305
"1890",-0.00643001588811876,-0.0133332273319198,-0.00330832670242698,-0.00453231864625436,0.0112116710614041,0.00457758478854164,0.00307144892963618,-0.00904615482896631,0.000393662424665209,-0.00267273931650935
"1891",0.00448442150029815,0.00395004217394779,0.00663877645005262,0.00569098266202372,0.000798891256444945,0.000193588325812399,0.00222722575297385,0.00890023940548268,0.00605962068151422,-0.00689125536772417
"1892",-0.00395691846923907,-0.0124250013793641,-0.0173124132467447,-0.00543233043319746,0.000265237570493015,0.00213240121390013,0.00319449357669055,0.000678752549222006,0.00547557119760866,0.00154199887714679
"1893",0.00137537323352244,-0.00062894568230043,0.00167788195281715,-0.00113787441312974,0.00637998777071003,0.00164447680416124,0.000692234628943744,-0.000451966127483439,0.00186716985428803,-0.00885304054897218
"1894",0.00503510556784259,0.00692399995702764,0.0117254072017992,0.00774677541212232,-0.00431434026718625,-0.00222099339004767,0.00456559508628573,0.00407047022237705,-0.02376143829602,0.00388352215418641
"1895",-0.00187250262869088,-0.00416759085923279,0.0033110649022825,-0.000678498375784597,-0.00203397657284698,-0.000871172975120738,-0.000275333353069618,-0.00045046167350915,-0.00946549467494828,-0.00928428552675742
"1896",0.00370116069219661,0.00795143004416121,0.00165010312461344,0.00248873402945815,0.00531654117052316,0.00145294449050959,0.00371934704069088,0.00743562534759445,0.00353330124093221,0.00156178810632168
"1897",-0.0113660143056721,-0.0153622471794441,-0.00658972096016563,-0.0187317858024679,0.0126034644351471,0.0058040107789068,-0.0059015410668295,-0.00849912184379198,0.0169640312317834,0.00233922971859379
"1898",0.0102192356498054,0.00780110136458978,0.00497512084844276,0.0156393866700477,-0.00322049207413189,-0.00201919883064305,0.00883598176141542,0.00924851782663927,-0.00755369447017684,-0.00661216291621969
"1899",-0.00187110504991306,-0.00460270338745894,-0.00165010312461344,0.00339685231701847,0.00497767403531868,0.000288581523612663,-0.00287401103832619,-0.00223513118886354,0.00166494097355763,0.00469848805988504
"1900",0.00435783175959314,0.0048340032363694,0.00330566093065765,0.0092530269944131,0.00208529644153588,0.00125259759419083,0.00425451547519828,0.00403239088171237,-0.00474907407785574,-0.00428688944394529
"1901",0.00221977934950601,0.00104600018468748,0.00082382879548093,0.000894417028029615,-0.0013007042423806,-0.0000966708878969991,0.00218713938827553,0.00401570360614412,-0.000954310497126021,0.00273980957205633
"1902",0.0000505949242759485,0.00522354548353987,-0.00493826790301011,0.00446824334374551,-0.00746656879615892,-0.00404147879085226,-0.00259125941611504,-0.00177754724656864,-0.010109894679751,-0.00117094414663099
"1903",-0.00468150300048176,-0.00706720997516019,0.00330848650622451,-0.00400360975153968,0.011808763896151,0.00386512680153639,-0.00560542009956344,-0.00823682804401638,0.011580241440776,0.00390772288067054
"1904",0.000404282020254332,-0.00167476828993551,0.0057709181847474,0.00692274758661027,-0.00138289139478665,-0.00115486643150586,0.00604928434762275,0.00157133884875305,-0.00166944111877387,-0.0019462560111887
"1905",-0.00429706679931485,-0.00293546920871357,-0.00245915011183928,-0.00598797266322837,0.00363570708553373,0.00134843336988677,-0.00464622691815098,-0.0011203855389984,-0.00302599931476344,-0.00312016237850077
"1906",0.000152204984740001,-0.002102965313448,0.000821797957220927,-0.00490861405770548,-0.0138875161803136,-0.00702419085159545,-0.00096134550891902,-0.000224433664764989,-0.00295523170020529,-0.00430358089483418
"1907",-0.0197481813718832,-0.0195996997104635,-0.0147783360626681,-0.0174887464075032,-0.00297429910398128,-0.000290782289845359,-0.0144312624629143,-0.0130166387191458,-0.0115357123842711,-0.0051080660694437
"1908",-0.00305550397198395,-0.00795352319120701,-0.000833348015211843,0.00547709131786411,0.00774112932930882,0.00588578948693286,-0.00195213985720288,-0.00250079301392514,0.0080233244835346,-0.00789890821798944
"1909",0.00722063364566772,0.00476687837754586,0.00166817820474585,0.00930552873583079,-0.00261850440214983,0.000578829231295153,0.00600812432008269,0.00364713680251461,-0.0031355443753549,0.00756371398691158
"1910",-0.00969609351870815,-0.0116451092276776,-0.0158202430627291,-0.0152913196476985,0.00323787279067589,0.000482302899393661,-0.00888849066295239,-0.00885766355420681,-0.000967779675260627,-0.00474118489242559
"1911",0.000312525681183562,-0.00218230300063615,-0.00507613810192864,-0.00685086979927518,0.000610983468424253,0.000868657253317417,0.00182133421160491,-0.00779108774231496,0.0145313228094457,0.00635168079479187
"1912",-0.00541476897515647,-0.0113711875815454,-0.00340132653706415,-0.00390897364742437,0.00932838429876925,0.00452905022914485,0.00153872962744983,-0.00461889534193827,0.00405826377111906,0.00197235968110299
"1913",0.0115687111299798,0.00906903523083291,0.00170651462145122,0.00900268073569443,-0.00215912499300353,-0.000863494076007609,0.00754202510872615,0.00556839424054556,0.0000792677127912089,-0.00472426408615978
"1914",0.00289808767491384,0.00197271146984512,0.00936955853143528,0.0128119716818922,-0.0000867502889010385,-0.000479894800374581,0.00554478529819069,0.0108447601937882,-0.00182267213213938,0.00158217528215698
"1915",-0.00139304197880541,-0.000437373180446676,-0.00168779351044523,0.0011292099574538,-0.00649296011949907,-0.0014412721718331,-0.0028950091265606,-0.000685075689544901,0.00023816291075085,-0.00631915096339819
"1916",0.00676881075107327,0.00415839380499072,0.00845323486717686,0.00541537914404144,0.00653539417323112,0.00327096784466496,0.0124429430909261,0.00799487833767776,0.00166679104161904,-0.000794901731337117
"1917",0.00472190946173545,0.00566705618657903,0.00167629025140603,0.00157071403157749,0.00805123995855261,0.0020139004773283,-0.000273261093925892,0.00702440655821746,0.000871640274286101,-0.011933134359741
"1918",-0.000204382470188946,-0.00130053321887669,0.00167366977735872,-0.00268873984796503,0.0109067828144016,0.00401896320246475,0.000956114252252727,0.0036001407279771,-0.00657109502923114,0.00402575128422056
"1919",0.00837948535336097,0.00781243489380379,0.00334183880638261,0.00966072963624987,-0.0099400853375613,-0.0031453853914567,0.0092796937948858,0.00470870217038155,-0.00414411848555662,-0.00842021728674447
"1920",0.00521870324016338,0.00193808331805867,0.000832562123295411,0.00467286279217327,-0.00308846812722918,-0.00105172701477896,0.000811093808611885,0.00490986589568609,-0.00224070904481988,0.00202189146360765
"1921",0.00267157824176834,-0.00429835960219038,-0.00582372971927625,-0.0019930745917921,-0.00163546072216592,-0.00296714699552625,0.00486347244181373,-0.00621832472781969,-0.00368943695861412,0.00282482003879458
"1922",0.0029157710770491,0.00561180819979312,0.00502110171835235,-0.00421703096663106,0.00560355554956993,0.00211198901210885,-0.000941006634822217,0.00335216352851986,-0.0107873449461653,0.00241449533829319
"1923",-0.00155396804155539,-0.00515137952089539,-0.00749388643207327,-0.00267407618834303,0.00557317770130217,0.0000956635108981807,-0.00672865231385011,-0.00178175124713997,0.00252282721002994,-0.00160580016755862
"1924",0.00507045839948672,0.0101404147117317,0.00335585652442183,0.0073742574514537,0.00375105742360793,0.000766430427000309,-0.000406439644868417,0.00401570360614412,-0.00365292631458847,0.00160838290910359
"1925",0.000649585390639196,0.00170867416802767,-0.00501690247234454,0.00598930033267608,-0.00322764116956376,-0.000191151445574023,0,-0.00133275429430091,0.00496985505898406,0.000401439712543361
"1926",-0.000399269944933667,0.00405138749205491,-0.00420166215635942,0.0050716757263507,0.00852174350913137,0.00277595576934009,0.00162641962088683,0.00311515828026709,-0.000243194166894112,0.00160511449347278
"1927",-0.000549738606916983,-0.00594619455051126,-0.00253159709976403,-0.00987275031880586,0.00523857335756706,0.00133627499470657,-0.000946930622074293,-0.00510232150350287,0.00551410963347387,0.000801271114856617
"1928",0.00284838377464713,-0.000213750150684811,-0.00169198376573565,-0.00155087584724245,0.00067254847629572,0.0000954433574440472,0.0050114819431335,-0.00267549923302568,-0.00112902419354843,0.00200165638693472
"1929",-0.000498490474160618,-0.000854778194150363,0.0101693892430028,-0.00155366857260508,-0.0172506092070147,-0.00638856349748784,0.000538730411072885,-0.00268276924397703,-0.0178427174403138,-0.0143828316073027
"1930",-0.00054832203483024,0.00940974231934266,0.000839033595195993,0.013114009721503,0.00556832216281555,0.00144186140595259,0.000269662740800092,0.0100872768968747,0.00411015200805331,0.00405353459188329
"1931",-0.00144630653196964,-0.00508467898542864,-0.0033530432085237,-0.00263280086639717,-0.0121824609693276,-0.00355081934866686,-0.00188536048470256,-0.00754550270816667,-0.00548505107678998,-0.00403716978450852
"1932",0.00449537884780971,0.00212948795018186,-0.00420510314448175,0.00857891115731668,-0.00189769060985134,0.000288851318589245,0.00944430202370894,0.00178913924068813,0.00477440719193911,-0.0016213804612808
"1933",-0.00258564089515245,-0.0131746791104084,-0.000844702684283161,-0.011777460437178,0.000432169360928825,-0.00105902101302602,-0.00173763191977094,-0.0111606255613018,-0.0108962397328566,-0.00487208260272087
"1934",-0.00633136829311776,-0.000645874643202093,-0.00845314154376242,-0.0123591692201792,-0.000777005905659434,-0.00231317659493036,-0.00535541335656575,-0.00835226040537485,0.00115961232933959,-0.00815990734283745
"1935",0.00376276304611189,0.00409388113083309,0.0110827964510167,-0.00424575492776891,-0.0063100229960128,-0.00251239668561087,-0.0138644170822897,0.000455249813114733,-0.0050467525842619,-0.00699312305008326
"1936",0.00114966117732029,-0.00450641296740861,-0.00252955558192003,-0.00673251121136564,-0.00330588604900162,-0.0012588731274259,0.00122838635051847,-0.00750859611322197,-0.00656910848878922,-0.0049708498179174
"1937",-0.00584145510520295,-0.000646775118960941,-0.00338101397662771,-0.0106191913111048,-0.0104728355706812,-0.00378159737056438,-0.0287663149384199,-0.00320955475768003,-0.00912366276786081,-0.00791018072039307
"1938",-0.000753235439339583,0.000431470993706107,0.000848097593119324,-0.00502396592075127,0.00149974294796595,0.00184912201533671,-0.00407091898053114,-0.00850924029643496,0.00219633389583551,0.00125898658360835
"1939",0.00753838044394262,0.00366534672922247,0.00169485142683512,0.0130823595181617,-0.0040515451099985,-0.000291318107441318,0.00747034145399628,-0.00139220700037079,0.00160150877951359,0.00922045596687138
"1940",0.00134697148308871,-0.00386690507582399,-0.00846019903576078,-0.00928858584736569,-0.00256396626070687,-0.00252720914129567,-0.00069949782929557,-0.00627161514852337,-0.0108558527163871,-0.00415285260395082
"1941",0.00532988509792753,0.00927330998280995,0.00597280117507992,0.00137203807287034,0.00319129339471558,-0.000681506263483178,-0.0072800395174647,0.00467478008265809,0.0020418410580072,-0.00959132395730922
"1942",-0.000901006675741223,-0.0049144681111537,0.00169619518623843,-0.00753589622728934,0.0127251191461299,0.00380249552429501,0.000563993256888162,-0.00503663256407916,-0.00585840555152328,-0.00294732818754173
"1943",-0.00772293727396367,-0.00365049431041198,-0.000846661489975475,-0.0151864730820531,0.00122197356552989,0.00213658909645442,-0.00887916469109262,-0.00329635082906143,-0.00204968834399821,-0.00844604763001489
"1944",-0.00572435884134215,-0.0129311063791343,-0.00169503854816311,-0.00560748524492705,0.00618770249249811,0.00213227318234521,-0.00568823992046219,-0.00685113531231718,0.00641848534734257,0
"1945",0.00782786040185357,0.00458512820327051,0.00594228629992566,0.0143326036156928,-0.00554338295423407,-0.00280481926141141,-0.00101039269057224,0.00404410485261297,-0.00467682831083038,0.00425901741067269
"1946",-0.0161353952438306,-0.0163007096315814,-0.00253159709976403,-0.0217744228670216,0.0118455137115743,0.00484982312063309,-0.00491190295369659,-0.0156363340030403,0.00290470731555637,-0.00212041208275215
"1947",0.00794547665620504,0.0041979806076069,0.00761434725643406,0.0044991139688908,-0.00146318532058243,-0.00212374779780322,0.0110336642492637,0.00890469953768691,-0.00281115088858641,-0.0016999779678657
"1948",-0.00181912744402046,-0.00748082521714721,-0.00587751663566827,-0.0202730904537596,0.00801698396875139,0.00319245584335315,-0.000287150593582419,-0.0102574517752779,-0.000256270293119143,0.00595994531177846
"1949",-0.0026322582874907,-0.000664785952822267,-0.00591217283331169,0,-0.00564437705180543,-0.000867729803983974,-0.00603265002513642,-0.00192816320094313,-0.00700675046575028,-0.017350806458111
"1950",-0.0135521475698703,-0.0126444098208419,-0.0161426679298911,-0.0204523965221929,0.0193909883797474,0.00840122560049905,0.00057797082924016,-0.0074863603545936,0.00481884523551201,-0.0034453030602557
"1951",0.000154506451746528,-0.0112333825902222,-0.018998415027047,0.00540417729079357,-0.0087115211746821,-0.00297172950895297,-0.00158868706210924,-0.0065687487146977,-0.000256906746345154,-0.00388940490539325
"1952",0.0110095153618641,-0.00431713346539098,0.0123239669742758,0.0085508194527093,0.00426621650546388,-0.000288624294769835,0.0067986548266854,-0.000734895702450444,-0.0182456487621321,-0.00954442786635024
"1953",-0.00117086714949788,0.00821546634798209,-0.00260874167022973,0.0130816476724711,0.000594683516779826,0.0016352877432162,0.00129313630140282,0.00171557006073741,0.0123898262595776,0.0127025911314935
"1954",-0.0154359864062856,-0.0212765603557168,-0.00610288875602294,-0.00884765734460735,0.0135010011811756,0.00585818947505801,-0.00588295694379293,-0.00831928317760122,0.00284410930659407,-0.00389276939652727
"1955",0.0174892145859415,0.0191949776847142,0.00614036270654261,0.0149577285695417,0.000251319821568785,0.00353211323233338,0.0190529458804605,0.0148039425174482,0.00953936052303739,-0.00390789288984161
"1956",-0.0198331700791865,-0.0297254391057566,-0.0252833378359445,-0.0156879393396611,-0.00435560985562544,-0.0017123877438463,-0.0012749794337128,-0.0133724119867671,0.00144716096495134,-0.011769807888793
"1957",-0.0114142500477286,-0.0137979718784673,-0.0143112268451656,-0.0217340732323151,0.00992685271561689,0.00390748817862274,-0.00141800236754075,-0.0056674062365234,-0.000425051006673338,-0.00352893522585584
"1958",-0.0164268975450595,-0.000236960144517684,-0.00907436979925347,0.0101209997910858,0.00608052213351584,0.00522129299605134,-0.00170415076223185,-0.00322160553782214,0.0079088445585116,0
"1959",0.00154731022265397,0.000711554948425785,0.00641016697532604,0.0058652249994724,0.00654080009022828,0.00198280631751935,0.0150802372291698,0.00273464545452806,0.00059060919483489,-0.0150509295657192
"1960",-0.00676639032757131,-0.0106658754323399,-0.00545932891499223,-0.0126337141865459,0.00789700970098073,0.00565515713527343,-0.00700778593150908,-0.00223161318867771,0.00337298265867214,-0.0125843292251807
"1961",-0.000857887548904035,-0.0103019467880785,-0.00365969112355402,-0.00910432770019698,-0.00636606770368431,-0.00271757744261913,0.00268206677852589,0.00447283437968071,0.00193296078549388,0.0100137531760711
"1962",0.0118106256751929,0.022028431614425,0.00459124599591498,0.0111745717836016,-0.0055851860999796,-0.00291369692691434,0.00506735921204648,0.00890698673417778,-0.00192923165635606,0.00360527101475738
"1963",0.00970971316886882,0.00450005450281532,0.0201097416087974,0.00294703034853505,0.00363451782392232,0.00141385264692362,0.0142855829892823,0.00882774805958952,0.00680733686540624,-0.00718459324177123
"1964",0.019811009636477,0.0150908630447992,-0.0017923193732039,0.00416261680427921,-0.00798304523710403,-0.00272900287800171,0.00952784033843646,0.0109380428085741,0.00183634386052556,0.00814114085177753
"1965",-0.00711076487624351,-0.0111499271797214,0.000897682059160632,-0.00658350643739647,0.00107825743280565,-0.000283258202990799,-0.000410162513256762,-0.00769407593866367,-0.00566573085316779,-0.011215776547182
"1966",0.0116247800312019,0.0136247400939751,0.00627813864170013,-0.000245795352984968,-0.00886675956290139,-0.00415361046522189,0.00752601038115541,0.00993458443744522,-0.00687111636906701,0.0117966179513764
"1967",0.00769512815166462,0.00463516674539299,0.00356529763845637,0.00712036389826043,0.00100327174393167,0.000853146500034985,0.000407520855211452,0.00239912656490371,-0.00143434866944858,-0.00627794142929505
"1968",-0.00137449247612964,-0.00553628578577792,0.00177586225491777,-0.0078012232016248,0.00183764423875776,0.00104188467667976,0.00597312100647507,0.00191468139568474,-0.00245035914576019,-0.00270768346460881
"1969",0.0114702245573752,0.0153096813861473,0.00531934142992463,0.0201472154229545,-0.00625321123965428,-0.00245996738094278,0.00323872841473749,0.0102728089519206,0.000338810779922261,0.0081448253341041
"1970",-0.00151212071051454,-0.0105096183866737,0.00529090368544405,0.00144517931296662,0.00226535729621857,-0.00331983575560602,-0.00739831845785743,-0.00638510573678353,-0.0143098562965259,0.0116697308327325
"1971",0.00641074866143043,0.00600311885017191,0.0078948765643525,0.00937952734353309,0.00083704126996631,0.00104675697166545,0.00853766928632615,0.00975766032359582,-0.0104802161161337,-0.00842948025412049
"1972",0.0114354117148749,0.0119351097722056,0.0496082172985688,0.00428880485277294,-0.00259302446859955,-0.00161632586158766,0.0075249709105607,0.0254535415487167,-0.0219636943838234,-0.00134235562090357
"1973",0.00054541209531056,-0.0131552380292109,0.00663343343551359,-0.00830362484656633,0.000000145506561022302,-0.000371744070653768,0.00773541851921378,-0.000919212938876091,-0.00452691267435068,-0.00896049769793583
"1974",-0.00346915314508711,-0.00229814915447291,-0.0263589975161229,0.000956677171995324,0.00311013438498997,-0.0000954387299310078,0.00119095409233871,-0.00897167498105034,0.000624155138222893,-0.0144666273901938
"1975",0.00631620448754067,0.00691084718538404,-0.00507613810192864,-0.00884290703001622,-0.00142445367882149,0.00028584183515945,0,-0.00789205999746312,-0.0216538939435582,0.0027524450020886
"1976",0.00400295342445078,-0.00388916103896275,-0.0127552326809737,-0.0122981369774877,-0.00646191671865359,-0.00305244430307428,-0.00422987099817185,-0.0138047356795331,0.000819710348668234,0.000914806340723828
"1977",0.000935088026441599,0.000229504063522956,-0.0034451053695832,0.00634748980717625,0.0114873550356647,0.00641144651368752,-0.000796714988695379,-0.00450740184159026,0.0281216243571611,0.00457041564431049
"1978",0.00314752892188919,0.00459256604667901,0.00777870751856002,0.00266888108981767,-0.00918547623144472,-0.00408877912636274,0.0045171645264126,0.00762622770692656,-0.0222183055482137,-0.00955414996961046
"1979",0.000980579270571047,0.00731410692745627,0.00600325192321027,-0.000967863166050797,0.000673976989625125,0.0000954827466062014,-0.00251283731023955,0.00614935041139897,0.0143038386230658,0.0050528032285897
"1980",-0.00107726720999901,-0.0115723628757401,-0.00511499202506038,-0.00193762958632515,-0.000842433511151097,-0.000381915878452155,-0.00517105661539929,-0.00376107748513255,-0.00481971612977761,-0.00319922509623971
"1981",0.00112730865722122,0.00367296413410689,0.00856903687474753,-0.00266930461113801,0.00236075790434565,0.00162378932980656,0.00399848505588341,0.00283145744469482,0.00152464573991029,-0.0183402430648723
"1982",0.000245208245272188,-0.000914887486839877,0,0.00827245613867289,0.00487749770619295,0.00209740001766323,-0.00610628075541964,0.007058770137363,0.0250739057056308,0.0107426411771041
"1983",0.000636308167407451,0.00228939458370814,-0.0161426679298911,-0.010617652855996,-0.00251102279711457,-0.00114154901247099,0.00373960258557804,-0.00420568471098648,-0.00366906609881124,-0.00415900323180507
"1984",0.00577376628975679,0.0139332914814712,0.0138169056043365,0.00536572831890147,0.00276901052351608,0.00114285363591038,0.00479060668075282,0.00375408243366948,0.00876808394297024,-0.00510438663375412
"1985",-0.00160534261118073,0.000225509955279257,-0.0059626258668557,-0.000484999391967667,-0.00635885023845062,-0.00266431677554069,-0.00622471815671488,-0.0021035855032594,-0.0119078919102679,-0.00513052706809547
"1986",0.0017541583634304,-0.00427942536382431,-0.0102827922180972,-0.001699035096146,0.00522096751592649,0.00181284132433057,0.00279854523044221,-0.00960406461843266,0.0103800228712174,0.00843884767950143
"1987",0.00535084289888288,0.00814288615393255,0.00779208253757169,0.0318504071461472,0.00603089459292816,0.00200029100564603,0.00730928322788937,0.00946044937102108,0.00461429562411375,0.0106925542322909
"1988",0.00280625482623953,0.00830139522485496,0.00171843330820365,-0.00824720895009223,0.000832391257866272,0.00114024653996481,0.00290227672272692,0.00164013031043941,-0.00242653611601129,-0.00873962635098224
"1989",-0.000723981113740946,0.00356057260429932,0.00257292031841283,-0.00641468818865087,0.00831938968088664,0.00246826189731286,0.00276222042227392,0.00233920669682197,0.00234554771657081,-0.00464030806755011
"1990",0.00255909292293088,0.00421279429609123,-0.00256631738826107,0.0126731423413704,0.00272307928974347,0.00170424711481476,0.00747765947172141,0.00210056463584052,-0.00190668231686641,-0.00233111440108369
"1991",-0.00211880141602983,-0.00684489993077086,-0.003430520972869,-0.0200707725596551,0.00789922547028366,0.00387602842093049,0.00286435627172454,0.000465675427002932,-0.0264849157177869,-0.0457943004701402
"1992",-0.00695008911924722,-0.00111152138036397,0.00516350681322431,-0.017108269721155,-0.00583422048996485,-0.00245237082403527,-0.00363547348779247,-0.000232681506243004,0.039871563287204,0.0205680919931677
"1993",0.00646393942946211,0.00022240392287709,0.00856153422095862,-0.000245154939674141,-0.00971200171404929,-0.0044447048596189,0.0035186914798131,0.00651899056959704,-0.0123520584602493,-0.0211132512505544
"1994",0.00386308552540604,-0.00177973245991547,-0.000848817711827543,0.00269733733879529,0.00390657691944885,0.00038016580099387,-0.000909299194186475,-0.000231006467610761,0.0103352701957204,-0.00588237341865872
"1995",-0.00110632967474888,-0.00401268678836642,-0.00254880404454405,0.00171188784848031,0.00836133422377472,0.00351320670337985,0.00155977785263239,-0.0115689350087295,-0.00386834859677898,-0.00295853949162506
"1996",0.00163728455684553,0.00492368540947274,0.000851709656438215,-0.00195324049710921,-0.00582912434340066,-0.00558257153346953,-0.00519062615465693,-0.00304316798334092,-0.012512918860362,-0.00247276535029672
"1997",-0.00668264231262183,-0.0075723567706264,-0.0161701452955415,-0.0146770004066017,0.0122222792611757,0.00333014734030468,0.00443494756520435,-0.0150271645268342,0.01179759678406,-0.0173525206683872
"1998",-0.000677677779427621,-0.00875202656132246,0.0051903069987751,-0.0094335256581819,0.0051401205911521,0.0036980011997485,0.00337702341176072,-0.00142999598049365,0.0208153655278578,0.0070634753146015
"1999",-0.0160311861604778,-0.0115462688620904,-0.0154908054695814,-0.0147873767954564,0.0073049496930655,0.00453566966811136,-0.00233012918485298,-0.0057291889447566,-0.00194604447168056,-0.0155310053935875
"2000",0.00506956133124126,-0.00366484993245508,0.00262252088239556,-0.00839487787163651,0.00410978800187545,-0.00169312414040934,0.000908213668329827,0.00432161015244703,-0.00228888608247602,-0.00916028487234122
"2001",-0.0161612914915008,-0.0236780160371198,-0.0095902125084002,-0.0164187311919691,0.0135623632293331,0.00819640940518496,-0.0090734249084734,-0.00812815951179824,-0.00237911458273243,-0.00821792272696698
"2002",-0.0068693568146837,-0.0174241599497803,-0.0193663448847241,-0.0143453579749814,-0.00205853555681124,-0.0036438527040239,-0.0117722899014293,-0.0110869961852751,-0.0257218711959162,-0.0160538006646467
"2003",-0.00801971131831225,0.0119818210261655,0.000897682059160632,-0.00158770132459463,0.0123770291885255,0.00506459746760379,-0.00463281631626822,0.000974840123615373,0.00489551538504673,-0.00578939496770725
"2004",0.0196048986668478,0.0108927894289073,0.0167812677476469,0.022986962522956,-0.00901275654318989,-0.00690576516976393,0.0223405605298945,0.00998316387807985,-0.00591561563938092,0.00582310723543245
"2005",0.0247290143658576,0.0210821830052867,0.0159715102947253,0.0136662412848372,-0.0177933460350466,-0.00563802112817002,0.00897512269568379,0.00867884129364382,0.00770110285379633,-0.00315774346202635
"2006",0.0042545582350364,-0.00145481326348107,0.00524023161735099,0.00700032798751882,0.0134455905392292,0.00368555645992208,0.00206252208766888,0.00320398783677045,-0.00330008678592986,0.014783378020544
"2007",0.0046000725727926,0.00439397108370221,-0.0026065169622409,0.0139032110729185,0.00135101906177426,0,0.016467358668556,0.00816533964232069,-0.0193429821210155,-0.0182101106723288
"2008",0.00134960550243091,-0.00368402162166714,0.00174237046414993,-0.00914173714217836,-0.0198351163001012,-0.00828556531482161,-0.00506270933511144,-0.00119109410964247,0.0016880941353683,0.0100688091195851
"2009",0.0000961850501668415,0.00670216990315242,-0.00173933988969899,0.00230671648663994,0.00544298677066535,0.000722674950670799,-0.00411289472333443,0.00166963050524305,0.000266090123578033,-0.0131163498056155
"2010",0.00322474598992617,0.00114782080415687,0.00696864536199371,0.00792615107076888,0.00371117027911483,0.00133027527795293,0.00387193392114438,0.00428555985254087,0.0182673144879129,-0.00106324961847593
"2011",0.00134340591149829,-0.00802577674385496,-0.010380664721692,-0.00608830753129008,0.00747508402292807,0.00341527019498877,0.00437115816425959,-0.003793274039531,-0.010101924408222,-0.00957959621759008
"2012",-0.00536608045339848,-0.00970872253785471,-0.0122377281913792,0.00204179967633,0.00271268057446505,0.00113519177045118,-0.00102428544944289,-0.00309362514193323,0.0134600072747426,-0.00107467628639846
"2013",-0.00992283895123325,-0.00723631444683215,-0.00530979239982809,0.000764378862349702,0.00190969877612468,0.00113350436722182,-0.0153764459778245,-0.00763887327641077,-0.0140624569634321,-0.00753093793412274
"2014",-0.000535427741436667,-0.00493768360138735,0.00177937893267588,-0.0132349292652906,0.0111181911006659,0.00509486821688476,0.0123630063346567,-0.00192472927651,0.00440218340549059,-0.0119242345282613
"2015",-0.0180594801542838,-0.0300093745561554,-0.0115452853689315,-0.0177972190337414,0.0157084377171937,0.00610161895375505,0.00334285937574563,-0.0060256084099366,0.0150771473513824,-0.014262180473698
"2016",-0.00941889794425865,-0.0107186678953123,-0.0161724123854228,-0.0042020967506543,0.0180173544944739,0.00671757772430315,0.00730278288372666,-0.0033946369316924,0.01139896343526,-0.00946031160562877
"2017",0.0124611326218937,0.00935739009351133,0.0146116546453259,0.0216249296350519,-0.00197489751185609,-0.00018559048599498,0.0129735726293938,0.0167884993814513,-0.00589141890646971,-0.00617957602536812
"2018",0.0177450031356421,0.0153693759164921,0.0126013252997914,0.0170364489750403,-0.0132426370415136,-0.00407829147170624,0.00565047420173936,0.0107678669166,-0.00420852014085715,0.00395698354185292
"2019",-0.00801357453679274,-0.00624665633016341,-0.0106666131421108,-0.00329956729596548,0.0109522020554604,0.00493275971840901,0.00037475194503922,-0.000236501563094849,0.0113851990445886,-0.0016891660869599
"2020",-0.00783358993925376,0,-0.00359392967799532,-0.00814856794111163,0.00572200184397254,0.00351951369964287,0.00549187413447649,0.000946841463282722,0.0110864401997877,-0.0219966048061198
"2021",-0.00281275301824635,0.00435172230599434,0.0081154712312772,0.00872920280503742,0,0.000923059213694399,-0.00260711215123943,0.00828042562192088,-0.00337376861291772,-0.00403703159616031
"2022",-0.00603717617123245,-0.00192590442211416,-0.00178883013733744,-0.00559952443092659,0.00758599591314324,0.00461048462414415,0.00659604815251513,0.00375401650079854,-0.00160801450209835,0.0110017664138224
"2023",-0.00916042023959174,0.00603013919441375,0.0071683398209843,0.00230364805896288,0.0157354131433787,0.00853534472329698,0.001359964273699,0.00186990886703842,0.0251759004392991,-0.0137458120305932
"2024",0.0131140084857124,0.0141452535849231,0.00889672379222839,0.00842673492992851,-0.0127487866611863,-0.00737128526366104,0.00852013299528687,0.0177322472143784,0.0130642878606864,0.0191638030508074
"2025",0.00213281009831401,0.00732866500332419,0.00793665598630788,-0.00151942219880574,0.0132891391993246,0.00229206216161981,-0.00783551311539099,-0.00802396531516991,0.0137120473484831,-0.0136752043521947
"2026",0.00504795210407427,0.00774454534155367,0.0017498003254468,0.0220647590419611,-0.0115587273228831,-0.00475650490075907,-0.00148094571671398,0.00762652963222243,0.000241594208734153,0.00635480048784021
"2027",0.0148709290448139,0.00302742458570715,0.00436699147468222,0.0191064843590487,-0.00359855314089774,-0.00248171293901289,0.01952571554273,0.00366951344949062,0.00804958525196198,-0.00114808995632198
"2028",-0.0054828985999934,-0.00510781554772755,-0.00347848891319036,-0.00754802849357716,0.0139184908345082,0.00654198930620709,-0.00206083789489919,-0.000228162536320298,-0.00798530684376009,-0.00632181185090264
"2029",0.0023416537998584,0.0151689971996674,0.0113437967032428,0.000490572457125138,-0.0030422934414337,-0.00228880132075049,0.00983840057546104,0.00617161005327116,-0.00998152596035917,-0.0034702855386991
"2030",-0.0131904066210551,0.00137955581539972,0.00172557337283963,-0.00539473795320899,0.00156306700267916,0.0013765764388467,-0.00132298110988105,-0.00477082861059774,0.0114643794042504,0.00522343606937192
"2031",-0.0128244842921275,-0.0197427881295785,-0.00172260089859688,-0.0108478859312887,0.0163483155732311,0.00769670864915328,-0.00710588384779032,-0.00890204677591611,-0.00787784553251047,-0.0144341619889924
"2032",0.00924368598600789,0.017095783256863,0.00862796155625567,0,-0.00657991761366239,-0.00354623047507341,0.00169840414297018,0.00967304162213156,-0.0215523905615361,-0.00468652079010523
"2033",-0.0125748069204363,-0.0161177843698398,-0.0171085714191833,-0.0274179542610312,0.0177371437644025,0.00876013195642189,-0.0163480502316737,-0.0177918771427142,0.0222755461696662,0.0241318147701892
"2034",0.0123839793285003,0.010999259876896,0.010443907685892,0.0179393903595053,-0.00377576243294975,-0.00125064400601926,-0.0032004838436408,0.018810755026329,-0.00834345099255041,0.0137930332837239
"2035",0.0144613631176289,0.0217591303150735,-0.00172260089859688,0.0188822985175456,-0.0211663004520604,-0.00843683606988699,0.0092623046815834,0.00866215733932818,-0.0111909412055373,0.027777866916868
"2036",-0.00380795913304666,-0.0124602051029176,0.00517686215660551,-0.00494200140947287,0.00170875171923401,0.00164701993832117,-0.00293689731656577,-0.00949172499509388,0.00437834768166012,-0.0220628612013305
"2037",0.0100950563165061,0.0137645596818146,0.00858369068389164,0.00595979886024578,-0.0109791909013959,-0.00365376395429351,0.0104321818055175,0.0182520306259593,0.00172724951920977,0.0135363096736323
"2038",-0.00276539540869347,-0.0153882931395478,-0.00851063799977891,-0.0170326775576055,-0.0177016203449892,-0.0111844529404589,-0.0263571480949767,-0.0100825445916307,-0.0258642086717776,0.00278243448269144
"2039",-0.00447583309843191,-0.00390680601647742,-0.00944196319279633,-0.00150682995400431,-0.00160375662921808,-0.000463146799154712,-0.0047406550018213,-0.0140336162060201,0.00446728763037174,0.00998887909743806
"2040",0.0106532037107256,0.00945990753163373,0.0129980155235054,-0.00251512555461597,-0.00795379138264285,-0.00250478655520281,0.00350933327980818,0.00367325744661295,-0.00587393649196843,-0.0126373600584188
"2041",0.000580494543019228,-0.00617144969537564,0.0017110707235759,-0.00731208341090828,0.00184999976132683,-0.000371644794029069,-0.00212282687474707,-0.00251615515651882,-0.011817346063836,-0.00779065618397379
"2042",0.00961676846508031,0.0200091572190195,0.00683165462960056,0.0213361368558382,-0.00330872180702424,0.000371782965232548,0.0107646747491621,0.00986018884986617,0.00230627829503716,0.015142982519029
"2043",0.00411635700419666,0.00338223138493787,0.0118746237299321,0.0114397871967757,-0.0102685728413129,-0.00334748407322372,-0.00544902671733116,0.00681193957708115,0.00545429539643072,0.0110495723323076
"2044",0.00157324985893381,0.00247204993397987,-0.000838289552616778,-0.00221290833480858,-0.0150559338339986,-0.00709098130268104,-0.00286389999348258,-0.00270602778408391,-0.0166977534319948,0.000546553163430996
"2045",0.0000949441664259698,0.00403489508306776,0.0176171700155872,-0.000246262201608616,0.00593978066361767,0.00479212691135467,0.00849167568826514,0.00248745837256559,0.00284453059487055,-0.0120152404922721
"2046",-0.000713688091758868,-0.0017860800579419,0.00741985078914698,-0.00419031801281522,-0.00661350622735679,-0.00252493317639313,-0.0190689316374292,-0.00383477367904017,-0.00343814692928124,-0.00331676100198663
"2047",0.00600053463119243,0.0134198322045636,0.00900170161193881,0.00668300725761939,0.00293269571123655,-0.000562390180916084,0.00921486692837892,0.00543445229120332,-0.00569262539774673,-0.00388247916964912
"2048",-0.000141936473061821,-0.00441416296979091,-0.00567723851727209,-0.0100810858528179,0.0114586695603049,0.00459649050956368,0.00787967830368608,-0.00180156025034539,0.00130118842211302,-0.00668153796059567
"2049",0.00284087815498868,0.00620703994552607,0.00489392804119082,0.0144062200046851,0.0131261455455822,0.00663007023951545,-0.0188629261924157,0.0051894623034745,-0.00147273672355541,0.000560530484758237
"2050",-0.000849746168377741,0.000660900471314951,-0.00243496912933849,-0.00195880784798785,0.00431829318311983,0.000927500953125104,0.00215009985853865,0.00246903314169078,0.00381741273959024,0.0151261328873129
"2051",-0.00118155524704588,-0.00462350702168757,0.00895018430244687,0.000245509292087442,-0.0136677531568745,-0.00593111009940284,-0.00845673793546908,-0.0033586401096698,0.00319795168188297,-0.00827820277748603
"2052",-0.00340605388555471,0.00176969596710785,-0.00403200387587832,-0.000735873202563186,0.00840777814143179,0.00354268508363642,0.00712869083378065,-0.00292071219445356,0.000775428620660046,0.0111296806566363
"2053",0.00631337529624743,0.00154538450395614,0.00242903159293983,-0.00147280232479308,-0.0186263328384428,-0.0074438082463546,0.00391795330469247,0.00856236894259044,-0.00413226569792469,-0.0143092756386252
"2054",-0.00410391763020945,-0.00859790818168971,-0.0048465795018886,-0.00762069781011165,-0.00362599429291022,-0.00215649526868622,-0.00264365629921537,-0.00513854076202436,-0.0018153440525589,0.00614179367706202
"2055",-0.00421572379868862,-0.00378007189559282,-0.00487009415086281,-0.0108989424612065,0.000316678411104609,0.000751612388323775,-0.00833164089934946,-0.00763525463859704,-0.00311769288024866,-0.00887895921922588
"2056",0.00109404743604258,0.00334828383239105,0.00570965358251097,-0.00150270739794212,-0.00126527188019243,0.000563429381726266,0.00330979495565531,-0.00045271488234444,-0.000955616358651601,-0.00391931914536592
"2057",-0.0140643705816696,-0.0180202381329388,-0.00162201092772352,-0.0152998237827221,-0.0220920953087773,-0.010227323835386,-0.030448983001216,-0.0185646404204682,-0.0273043391304348,-0.0123666170244006
"2058",0.00414452664286546,0.0038514447612592,-0.00324933681977424,-0.00382038900211501,0.00923068811607641,0.00464556012718065,0.00889793121226057,-0.0129179130731153,0.000983372063442012,-0.00284572097699964
"2059",-0.0162220469003539,-0.0243736012175428,-0.0146700178441255,-0.0222451984262076,0.0131581596693253,0.00424587072722793,-0.00492842135082427,-0.0170600733274772,-0.0049120567570593,-0.0131278504276504
"2060",-0.00234170977092518,0.000693840728867468,0.00909833456138021,0.00758372895170401,0.00728490022575068,0.00178516706117415,0.00143368915060238,0.0028528779783028,-0.00601326523089696,0.00520530925471774
"2061",0.012713948633803,0.00809071098391101,0.0221313566920771,0.00622905861833267,-0.000707046357968033,0.000937879644817841,0.0165299383377511,0.0109058883929571,-0.000270871331828459,-0.00460298819676297
"2062",-0.00613209977962481,-0.00710851888856223,0.000801724232958767,-0.012122913761576,-0.00306834315213711,-0.00149929092277856,-0.00371304972305697,-0.00257988494799288,0.00144505056498345,-0.0202311155214705
"2063",0.0133604724594811,0.0145495212991478,0.00400657512476199,0.0120104040098399,0.00962724446924601,0.00347207964586782,0.0109243524804956,0.00940527028600946,-0.000631304129634969,-0.00118004618052503
"2064",-0.00297250156342999,-0.00409735271893918,0.00239415922983999,0.0116098352689851,0.00828532806774973,0.00205768853358768,-0.000890317329491741,-0.00652231946013015,-0.00541466483917807,-0.00708803408364778
"2065",0.0120215480207506,0.0237714760480221,0.0159236749201208,0.0244836631281273,0.019302404965436,0.0114788771378278,0.0197224795133171,0.0192260062619907,0.0195989839361128,0.0273645963994336
"2066",-0.00456114536958152,-0.0136190970295931,-0.0117556665402614,-0.0169281791877791,-0.00509537049866071,-0.00470538552243771,-0.00149711376194783,-0.00253031379261115,-0.000711951569494884,-0.0167920756911898
"2067",0.00882668575113743,0.0251245337297363,0.0158606240894079,0.0149407307345857,0.00527409596014627,0.00407849407522054,0.0242438622713426,0.0197232849749041,0.0113990470086467,0.0135453445761553
"2068",-0.00194861783412204,0.00507839386912567,0.00468354856579567,0.00299402513527025,-0.00121651975366821,0.00129307188165195,-0.00146421645524331,0.00136204239417292,0.00633971119133592,0.0116211714476675
"2069",-0.00561899911532293,-0.00175772126692186,-0.00233088957602501,0.00398009809595257,0.00966916363024484,0.00304284708195413,-0.00806467380252995,0.00702768289257572,0.00244989935733742,-0.00804142308010869
"2070",-0.0146538514199778,-0.0052814642363197,-0.00233627121046021,-0.0158575322919358,-0.00844534413430575,-0.0043211006395123,-0.0165174673487477,-0.00562815510085257,0.00139655232608882,0.00289521423429195
"2071",-0.00238147312668879,-0.00973462002946723,-0.0101484846111944,-0.0093151947823602,-0.0155895517733545,-0.00563149915099925,-0.00568222524626638,-0.00950858103682839,0.00653708690306587,0.0121247840176284
"2072",0.00228966019109977,0.00178735619696502,0.00394322838224292,0.00279560947732249,0.0124372975058609,0.00389991588374228,0.00342874352549716,0.00571446962333177,-0.00363703662182968,-0.0199657933908359
"2073",0.0121997728179213,0.00356846580023129,0.00392771885175724,0.0192600764548283,-0.00495953756084766,-0.0000929349601553886,0.0112643871204587,-0.00454552615656068,-0.011385346973498,0.0052385780379427
"2074",-0.0087393456920094,-0.0162223909796989,-0.0195616752858211,-0.00223789321725387,0.00214707043285212,0.00258998165677249,-0.00725905515564262,-0.0109588735374352,-0.000791173626373598,-0.011580737745951
"2075",-0.0035362547143859,0.00880949477522219,0.00399025808404541,0.0124598515469787,0.0131344577907631,0.00475923411838153,-0.00012628238303114,0.00738689869111675,0.0170683963727469,0.0181605695309341
"2076",0.00359736689385048,0.00806086194371347,0.00874401412662196,0.0150133509662291,-0.0105954193825923,-0.00285111353301026,0.00668272873096099,0.00801998134326731,-0.00276815748733827,-0.00517835431905656
"2077",0.00673309982430093,0.0093290944518083,0.0118203636307501,0.0128517513310433,-0.00558386955544843,0.00129115777778144,0.0100201177780386,0.00727451515979238,0.0122311156508599,0.0127241223596799
"2078",-0.00264615465172446,-0.00154041303352825,0.00467277747331374,-0.00502784568017167,0.00838449648870254,0.000829094016600029,-0.0162450182406491,0.00157982217772856,-0.0049704429690558,0.00513984965216796
"2079",0.0033770027705684,0.00110202962117567,0.00155040477698654,0.0209337201546813,0.000305405635316669,-0.000920269739904001,0.00277319779451468,0.00968854316538326,-0.00551201442156568,-0.0193180940344471
"2080",0.00442349888141136,0,0,0.0098985534144449,-0.0129646380966968,-0.00405381208200895,-0.0175988243517703,0.00290137877355301,-0.00692823238132634,0
"2081",0.00545697967166103,0.00330268277260681,0.00154800474303807,0.000700444784692777,0.00146821938318342,-0.000277354280131425,-0.000639983922063547,-0.000445093174625488,0.0113369061016291,0.0104287728250716
"2082",-0.00452296384120376,-0.00548598988262416,-0.00695505314556399,-0.00583059531913888,0.00138869540637598,0.00203555653383747,-0.00281687311956935,-0.0131342568854391,-0.0071570405522372,-0.00458721091733771
"2083",0.00191305908580675,0.00882609150868818,0.00700376470128039,0.00445707125339534,0.00708777810912076,0.00295498299881225,0.00205431011126178,0.0090233782975182,-0.00607952932151745,0.00460835039256935
"2084",0.00448722922750333,0.00503052802401416,0.00463683638439871,0.00700606357356559,-0.00084127731298933,0.000552583962616593,-0.00589401370649567,0.00268258153532042,0.00865080376353022,0.0200688264583102
"2085",-0.000285241580217255,0.00174088827940433,0.00230777044639363,0.00788502960325665,-0.0049766940234407,0.000735942897969855,0.0041243961238786,0.0031213908324188,-0.00346531231049119,0.0106800103349713
"2086",-0.0115034033836664,-0.0134692045023592,-0.00767461770413636,-0.0174873003140539,0.0114648659081171,0.00202268620641122,-0.00526286802098952,-0.0115579666313371,0.00495522042037044,-0.00222466379608099
"2087",0.00913692297183033,0.00110074747269251,0.00309363587932632,-0.000936727907797863,-0.00882465353362749,-0.00183520026825923,0.0012906157581849,-0.000674756786301689,-0.00761243092755071,-0.00445924791956631
"2088",-0.00119149265953622,0.00769927242978885,0.0154200509803997,0.00586005200605344,-0.00452850540512095,-0.00211429173078403,0.000773273096037919,-0.00224998694542666,0.0057531031576612,-0.00727885080943291
"2089",0.00491423824525805,0,0.00759326484951472,0.010720262629669,-0.0152659223334497,-0.0058038646411358,0.0029617199833416,0.00270629891828955,-0.0134338277023877,0.00338416449252255
"2090",0.00251628487734434,0.00545735166929484,-0.00075378404989479,0.00737844861047199,0.0043065851659001,0.0030580359339194,0.00179761211192786,0.00202442107324918,0.00729159259788115,0.01236644346353
"2091",0.00232057145084918,0.00434210781942901,0.00377081153217507,0.00366203384454189,0.0062367259697067,0.0035101122451151,0.00166642537725137,0.00606038540704579,-0.0140415222731023,-0.000555353763433186
"2092",-0.00415792057809983,0.0071336650823437,-0.0022539999253367,0.00387688114861562,0,-0.00156477014167999,-0.0026870232437145,0.00178504864305151,0.0201680578460488,0
"2093",0.00317889649483605,0.000429192922711596,0.0030120812369816,0.00159010517687674,-0.0137908243223016,-0.00461033966622182,-0.000256910413786726,0.00289523006805692,0.0086707706811624,0.00166675834314023
"2094",-0.00411464189753763,-0.00836732610612367,-0.00900888096510932,-0.012474452719755,-0.0122558674305132,-0.00370490450471506,-0.0196353629359834,-0.00644010923906957,-0.00704891245510331,0.00665542577805445
"2095",-0.0100204824514775,-0.00302888519676803,-0.0257576463027159,-0.0151581910979054,0.00174959594176793,-0.000279484258491669,-0.0116508569515892,-0.00916407744585057,-0.0176608169394716,0.00771362090786609
"2096",0.0108415585078776,0.00802941665633727,0.0124416656576911,0.00606325087772608,-0.0134612536719918,-0.00546661493407197,0.00529786652783359,0.00248123967549962,-0.00343702297138437,-0.0010934787598561
"2097",0.00284739021839364,-0.00172232641693915,0.00460828191806617,0.00579503450083285,-0.00943553014081433,-0.00206031743192425,0.00263525697217593,0.00607538822656006,0.0090201271839383,-0.000547337882276788
"2098",-0.0114520084094197,-0.0148801647055591,-0.0191131800286158,-0.0108319827198304,-0.00138395742626962,-0.00168896391190099,-0.0219451013435743,-0.0136432418663226,0.00280455745494401,0.00821473346996493
"2099",-0.0041168477320439,0.00678631743836444,-0.000779314134701559,-0.0123484096902768,-0.0171205628087628,-0.00488849872058117,-0.00268674222772358,-0.00680252310069007,-0.000524357638950534,0
"2100",0.00398964464258156,-0.00413161506182247,0.00155992948471528,-0.00141560853726708,0.0134376870850004,0.00425097473334968,0.0132023034808915,-0.00639280760151051,-0.00821968338387813,-0.0157523714176044
"2101",0.0131660449882609,0.0248910456962681,0.0233645925237485,0.0127569270041141,0.00270087361589888,0.00385672963946004,0.015290189318244,0.0238971037725901,0.00484925947538795,0.00551868825165203
"2102",-0.00477267283354454,-0.00447371407967145,-0.0159818147251406,-0.00956374531634241,-0.0243246763843087,-0.00983859962623923,-0.0145364335182672,-0.0089764691612737,-0.00386068260190675,-0.00439071958871129
"2103",-0.00299149906441032,-0.00385184411755113,0,-0.00329732025143992,0.00259331037171107,0.000756880716630937,0.00292362431524751,-0.00181172689154518,0.00854400606486383,0.01047394718828
"2104",0.000190627239138541,0.00644451306324867,0.00618725053898994,0.00189041247235577,-0.00801105400837931,-0.00132398213654505,-0.00834742459038162,0.0111159353438959,0.0179039563318777,0.00109120500779669
"2105",0.0104276624539168,0.016435507266118,0.00538041894624008,0.0099056376188642,0.00269233183924111,0.00340902701137602,0.0181720740812492,0.00964760835929424,0.00540537952624498,0.00599463697079994
"2106",0.00108384836478304,-0.00146996821217227,0.00458720599855567,0.00770678671368841,0.0200507506448329,0.00717180427794251,0.00826758290967922,0.00866672270801772,0.00298684929168802,-0.000541704379498187
"2107",0.00310672174492543,-0.00546800095877276,0.00837136113625192,-0.0101971548621798,-0.0167783080405877,-0.00674580994350626,-0.00299344298698379,-0.00837152798170682,-0.0000851016768919077,-0.00271010147902528
"2108",-0.000328465255402755,-0.00338319249250607,0.000754611304152775,0.00163906324432883,-0.0088666548523787,-0.00443385048490297,-0.00130561114765182,-0.000889042309883292,-0.0138699629136307,-0.0211955866319149
"2109",-0.000704211467629001,0.00297030207564397,0,-0.000701192335139544,0.00168811321783835,0.0021791078167972,-0.00209138418270882,-0.000444465104326053,0.00163951161998011,-0.00222107217221601
"2110",0.00291235456443006,0.00571191258716564,0.00377081153217507,-0.00350892686903936,0.0139861569393966,0.00595641169315009,-0.00458489644001869,0.000222466911058872,-0.00335975183735771,0.0122427460883201
"2111",-0.00238856313570546,-0.00946558843128054,-0.0022539999253367,0.00328640432791039,0.00041505358079319,-0.00225548061213099,0.000262775125013937,-0.00556091757759891,-0.000777975611064519,-0.010995183959485
"2112",-0.0107517593906556,-0.0205989716828993,-0.0128010870020421,-0.0159100578624916,0.0171097513888319,0.00621718534953164,-0.00605142667053449,-0.0138667516494407,-0.014619325512445,-0.0194552740661222
"2113",0.00949211884057966,0.0125759893870983,0.00686503166014663,0.000237569741526666,0.00228672262595886,-0.000561748865347322,0.00754485428008378,0.00249474600815924,-0.000175621098213563,-0.0136053739085655
"2114",-0.00112832136721552,0.000642361186398155,-0.00227294930095878,-0.0130734979443967,-0.00244422540466849,0.000936729370962341,-0.00065692204309209,-0.00610849910592204,0.00114143472773232,0.00517234311863457
"2115",-0.00621285917530789,-0.0113416669937974,-0.00911140532825805,-0.00963371896895659,0.00220508488247639,0.000561455651198361,-0.0107798213434477,-0.010243609128223,0.000701640081607779,0.0125786219037087
"2116",0.00203658854351629,-0.0069267116681756,0.00459766678518192,-0.0038912429800142,-0.0107477157772159,-0.004412476066322,0.00970137026704831,0.00184018619519399,-0.000876406676185937,-0.00225858023963132
"2117",-0.000992775662438716,0.00762868811093198,-0.00228838574334678,0.00390644390242634,-0.0139517063187559,-0.00696257477630557,-0.0081603021442197,-0.00114795332423157,0.00403507894736843,0.0118846210882944
"2118",0.00264963024221787,0.00865246077824411,0.00382255629571659,-0.00510699211497401,-0.016074795121095,-0.00852759937515846,-0.0120751204086312,-0.00459693495765356,-0.00716407484854154,-0.0128636462591393
"2119",-0.00844665975125103,-0.0113660913753573,-0.00685449194674193,-0.0151553741438544,0.013018844142064,0.00487370521145558,-0.000940627707875397,-0.0092356097231443,-0.00703980118831227,-0.00906514926579005
"2120",-0.0017132645827197,-0.014099881364222,-0.00613505748940291,-0.00446747525688651,-0.0121798966511384,-0.00722794562561879,-0.0120997973378734,-0.014681760823089,-0.0053172458460562,0.00457409782496465
"2121",-0.00614933852840194,-0.000439776898195188,-0.00540117770473147,-0.000249459535036745,-0.00110530947920839,0.00143734107700144,-0.00204120433431443,-0.00402115269649617,0.00294014616785709,0.000569144195399662
"2122",-0.000144158747924616,-0.0050628213489825,-0.01008516077969,-0.00598475326691716,-0.00791719225986176,-0.00325264661373703,-0.00722769669588563,0.00522474112848736,0.00222084036599446,0.015927265450697
"2123",0.0119933211509189,0.0250001374089068,0.016457589118495,0.0145509009524032,-0.00875224786600926,-0.00383855340842798,0.00714279188808775,0.0181905243223563,0.00850912072327614,0.0039193191453657
"2124",0.00322354387433244,0.00215810895991475,0.00462602587122962,-0.00494563869641684,0.0210351484410449,0.00789961874492739,0.00791032394161717,0.0025519553436244,-0.00457019691132188,-0.00892358463847098
"2125",-0.00765488143798276,-0.00969178155142347,-0.00537232925422215,0,0,-0.00057370199131479,-0.00189417603708353,-0.00485990087500454,-0.000264868439610377,-0.010129466925154
"2126",-0.00428544361392114,-0.0108743479161909,0.00308645379584593,-0.0111830294194445,0.00161097494966778,0.00239129639037339,-0.00515187299381137,-0.000697477704375227,0.00441579075114928,-0.00454797665417239
"2127",0.00545174591116226,0.000659592542260112,-0.00461543536576481,0.000251351507056574,0.00787192785981827,0.00381612778048157,0.00844918771051906,0.00023249729984598,-0.00360505573889769,0.00285547202898218
"2128",0.00161701278404447,-0.00131852250658471,-0.00850066527369675,0.00603040628956464,-0.00772614133111715,0.000570568978012664,0.00621615880329673,-0.00302466040572447,0.00467700317684439,0.00284745874768899
"2129",0.0103992734347453,0.0127612758825195,0.000779399674917247,0.00924051693191674,-0.00490948964043858,-0.000760163698208194,0.0138329588717931,0.00560090261532276,0.0129117437489985,0
"2130",-0.00443903847996807,-0.00391042163663313,0.000778856789350524,-0.00866131516689472,0.012843805232496,0.00532398457686112,-0.00649117595565019,-0.00359054688420024,-0.00173427852930974,-0.00908585572589227
"2131",0.00512308049707588,0.0233369764403284,0.0155643082626693,0.0144781454560401,-0.0204063474373001,-0.00841609450917824,-0.00986639586498761,0.0101271261706755,-0.0128561845155615,0.00343846653051139
"2132",0.000707936940804288,-0.00149189879780842,0.0114942615733715,0.00984296685423813,-0.00600103525827811,-0.00305157301438774,-0.00484808950386328,0.00373081212335546,-0.00659978886483448,0.0119930413004823
"2133",-0.00726287917923985,-0.00787782270091242,-0.0106061752419134,-0.0070665400187202,0.00862437300127827,0.00296517409229247,-0.00562483696386928,-0.00766574983207635,-0.00265748075699779,-0.00677197507159488
"2134",-0.00304057690223625,0,0.00200094895127445,-0.00343621660801496,-0.00350596255366298,-0.00247942083659625,-0.00947423208888276,0.000702457821972535,-0.00133221427594676,0.00113634815293406
"2135",-0.000190455103263543,0,0.00460824536493853,-0.00942703917383692,-0.0112408669236976,-0.00478081627270832,0.00485161325539685,0.000233706364646036,0.00106720026561358,0.00454040856141935
"2136",-0.0209702413849292,-0.0335599177383757,-0.0252293276893887,-0.0222890470382749,0.0264691711793792,0.0116246931628892,-0.0160020796013959,-0.0240877365798423,0.00453093469315813,-0.00451988643037415
"2137",0.00209317356493943,-0.0074896735778579,0.00470600310807434,0.014856686492843,-0.00693280013661679,-0.00275437978783455,-0.000420607032080134,0.00311530018104644,-0.00619082869019183,0.0215664003574805
"2138",0.00801557320702595,0.00548816611293446,0.00702550370490584,-0.000757276895381298,-0.0134980052872334,-0.00522638048857271,0.015287375199577,0.00334426851179082,-0.00347067713435945,-0.0122220558958132
"2139",-0.000915702148146291,-0.000227555667617341,0,0.00479897135631169,0.00328678377929981,0.00354764145781128,0.0022104071872695,-0.00214286224346794,-0.00196464541977193,-0.00168738161556348
"2140",-0.00284579215201186,-0.0245677349716027,-0.0069764903461319,-0.0279033805815906,0.0185344627353645,0.00706963058001464,0.00454827066109997,-0.00978257546353978,0.00268428771144791,-0.0326760730635546
"2141",0.00628861501337252,-0.000932660158998733,0.00234169250031036,-0.0149986344191603,0.00939456967922969,0.00265661786962679,0.0153680705713715,0.00192770770260053,-0.0116008925861304,-0.00582415211058229
"2142",-0.0167771654574497,-0.0147060623324706,-0.041277113883573,-0.0343921590137567,0.00863648791242011,0.00397352197550727,-0.00527043926885751,-0.0264551605399085,0.00297936072626648,-0.00468652079010523
"2143",0.00180889845130983,0.0175313452542929,0.0121851393413084,0.0193039335896199,-0.0197022423498231,-0.00697408712390013,-0.0047545443532282,0.00963423243949735,0.00243050688380619,0.0117715903659563
"2144",0.012591327925523,0.0419091852526328,0.0160512436389708,0.0253397400806632,-0.0158582383525389,-0.00692751496091748,0.0069612819024798,0.0200635076594387,0.00116735810733348,0.00465380499809842
"2145",0.0110372711003981,0.000670510026075766,0.0134282546171336,0.00676410669471195,-0.00310191318835717,-0.00267624004628275,0.0014912487038492,0.011513506151168,-0.00448470722907357,0.000579150118952709
"2146",0.0043381950479906,0.00848595749248315,0.00623526223221149,0.00180877159485271,0.00328479479212884,0.00316223693184936,0.00270685172636886,0.0075886414664883,-0.00225245521673045,-0.00347241290050826
"2147",-0.000332162998184948,-0.00465016463392798,-0.000774588654136932,-0.0113489354644414,0.0105968150263849,0.00382055837117101,0.000945116049820172,-0.00282415821184878,-0.00523743914100483,-0.0116142449742631
"2148",0.00802418897232204,0.00912121056879922,0.00387607250328981,0.0125228867586287,0.00690517602206664,-0.000380303251117819,0.00714763368243454,0.00991273794884528,-0.00363110008601675,-0.00470034876032666
"2149",0.000847932055312972,-0.00352723268709154,0.00231637725898737,-0.00128847965708123,0.00516504217129521,0.0000952118641133204,-0.00388343245185208,0.000467476408399392,-0.0101129735766586,-0.0053127963211177
"2150",0.000517864574542726,0.00309722139717716,0,-0.0064498949509455,-0.00421184174071132,-0.00199855444388564,0.00174785442499892,-0.00186918828344673,-0.0271514491090392,-0.0160238240596492
"2151",-0.0039513851646632,-0.00374954489879364,-0.00308151963533398,0.000259721032192406,0.00541382848488725,0.00276547250979076,-0.00362333602955445,-0.00397831585359998,-0.00312198684357579,0.00422195857957752
"2152",-0.00179473045024403,-0.00730565000555194,-0.00463675699066135,-0.0142784583605222,0.00622583531921372,0.00123637964702161,0.00282838025062881,-0.00258432343014736,-0.00540950919399696,-0.0144144029424824
"2153",-0.00562992913930527,-0.00289925648394773,-0.0007764775539576,-0.00974441460305298,0.012457927637757,0.00408519782065841,-0.00711787574262557,-0.0110722334831893,-0.0044847422380323,-0.00853139209343812
"2154",-0.0103720367211324,-0.0118540192592168,-0.00932384710298306,-0.0143618186766499,0.00247779091773892,0.000945719940694367,0.000270329056532015,-0.00261999714165895,0.00977663165385545,-0.00799018329028789
"2155",-0.00581738434187762,-0.00792222572319423,-0.00392167282514277,-0.0188882373332531,0.00535438971716395,0.00330818685268874,0.00216359673284017,-0.0028659455205895,-0.00465113440248954,-0.0192069322486307
"2156",0.0122832026447139,0.0134610549177325,0.00472459565792982,0.0101759842118663,-0.00729249855102032,-0.00282646493537764,0.00188917095020957,0.0124547492516616,0.0015258058218024,0.00821227311896955
"2157",0.00687906695014773,0.00225128234673089,0.00391853491639615,0.00980119979351812,-0.00371462937499356,-0.00141652871498654,0.00511792373066378,0,0.0014283089343452,0.00313291822478545
"2158",0.000237046235138649,-0.000224511003749872,0.00156114254033946,-0.00997548990683217,0.00770489902439087,0.00113464867901225,-0.00375188429283668,-0.00260205383224554,-0.00855758312365851,-0.00374779901424127
"2159",-0.00151778024232785,0.00629067759533952,0.0077942054521587,0.0108929637319131,0.00739978418147413,0.0058593690475468,0.00645606603847337,0.00308343118449916,0.00632974987042534,-0.013793109233514
"2160",-0.00337286521031255,0.000223183391360404,-0.00386701560442759,-0.0167023781202291,0.0105263497122803,0.00304826881843989,0.00494436550810007,-0.00425630330985316,-0.00791005432192893,-0.0165288315302095
"2161",-0.0019542277993484,-0.00267855688246499,-0.0015527219696605,0.00356143968703604,-0.00793214583821555,-0.00515924316451954,-0.00518598096229106,0.00403676162054611,0.00201729110503912,0.00581769849731795
"2162",0.00329537560405369,0.00671441581772791,0.00622073770422382,0.000273051013696346,-0.00750590548020769,-0.00386595185759619,-0.00427767601004048,0.00496717436646299,-0.00364296814577625,-0.00385605447913029
"2163",-0.00818776334985183,-0.00111153705525324,-0.00309121351933461,-0.00873333834375212,0.0088781688524866,0.0035023383753463,0,-0.00117694266281965,0.00442604637736932,-0.00064521886644664
"2164",-0.00191985563683705,-0.00400635118819781,0.00310079875035241,-0.00055082507439963,0.0131182094417468,0.00396193722457783,0.00349034484752986,-0.000942190366558626,0.00249068878715097,-0.0038734139922495
"2165",0.0125992669820036,0.0118437846350288,0.0146831903804423,0.0168043892638996,-0.0123853539738599,-0.00413436100810904,0.00013391815928121,0.00778260371318273,0.0102245482995786,0.0213869496870762
"2166",-0.00902338326983798,-0.0136926515694319,-0.0175171955821133,-0.021945527170855,0.0158794448753892,0.00660465946887423,0.00668788937468268,-0.0142752679097928,0.00510784141971388,-0.0133249515791739
"2167",0.00119837612677487,-0.00582180551762945,-0.0062013647238931,-0.0155121314609806,-0.00545093384906092,-0.000375211293437094,0.00146183838808955,-0.00261192343189698,0.0140221905887035,-0.00321539024234307
"2168",-0.0012446897647943,-0.00292790969153778,0.00780013558472614,-0.00168826630949626,-0.00322376824947834,-0.00262507636990483,0.00199000064322896,0.00166641918655763,-0.0082598515081207,-0.00451613365891079
"2169",0.00364229649226644,0.00158115622401045,0,0.00140912472966837,0.00234453103675603,-0.00103425349673258,0.00569389483031446,0.00617849155918604,-0.0000936084587908059,-0.00648092618506435
"2170",0.00558683865241649,-0.0036083994657059,0.00232207298760456,-0.0109766148308971,0.00451768699292421,0.0017883062694759,0.00750506081545033,-0.0002358114224561,0.00262048671259696,-0.00391384098282155
"2171",-0.00289676735475919,-0.00565889696587019,-0.00694978525142709,-0.0108141303035076,-0.00787021894348894,-0.00159724592010702,0.000783792174587017,-0.00519736207210519,-0.000186651736768018,-0.00523909389894606
"2172",-0.00790526204859865,-0.00956062708935468,-0.0108865510173918,-0.0123702778273158,0.00987528878443689,0.00611594026957851,-0.00548434842180534,-0.0047496176030023,0.0134441414112207,-0.0111914887418054
"2173",-0.0208813993183732,-0.0216043036348489,-0.0298740746775251,-0.0157297122051139,0.0100995745703374,0.00271207011974584,-0.00774649311363473,-0.017418389804244,0.0174113214902445,0.00266307934858157
"2174",-0.0301023695049794,-0.0216113315011982,-0.0340356874155635,-0.0307782449966864,0.00301540762111774,0.00401052116678224,-0.0195846645465282,-0.0206409083002371,0.006247690940824,-0.0166002437314864
"2175",-0.0421068572352798,-0.0268907403650331,-0.0352347493559865,-0.043664065287991,-0.000316412765666074,0.00167197476860426,-0.0467000571081171,-0.0453757449285994,-0.00539906430484294,-0.0249831944517125
"2176",-0.0117679328985676,0.00616823460473714,0.00608663294582934,0.0127713132356444,-0.0160651629519573,-0.00547155376811304,-0.0252017852514494,0.00701321261114485,-0.0123947798099592,0.00415521063827451
"2177",0.0383938486506736,0.0166746186529811,0.039758155772013,0.0331022442742623,-0.0193033959431833,-0.00615431474701567,0.0249817673421546,0.0201183932194857,-0.0136497429956122,-0.00620695348291322
"2178",0.0247350071635288,0.0108541480128057,0.0182875236997144,0.0442477717689365,0.00057405906026875,-0.000562916675905467,0.020121797286037,0.0199746815593678,0.000557304737759834,0.0360860590358638
"2179",0.000050227987950402,-0.00238624979150814,0.00489808526780733,-0.0128581554938907,0.00295084590399286,0.000187351177353579,-0.00111116692464241,-0.0101634722057422,0.00900393551460321,0.0261219592799926
"2180",-0.00807883901392081,-0.00454427197307561,-0.0154346650626789,0.00177612816816586,-0.00768235317751387,-0.00168939503115451,-0.019886012156765,-0.0120210201872664,0.00110398347113105,0.0241513737615482
"2181",-0.0298478545798284,-0.0285920378196035,-0.0453796633192231,-0.0387113111328014,0.00720548303764357,0.00449201677120503,-0.0190123808424344,-0.0263625830073452,0.00349197757765118,-0.0331421357263799
"2182",0.0189810216614221,0.0140983731490614,0.0181505388420207,0.0144481084537189,-0.00860440533814011,-0.00271880884373177,0.0107029137122265,0.0179639526698487,-0.00531130051221518,0.00856963182897941
"2183",0.000716421012260771,0.00146356178999585,0.00763988159923845,0.00393944162265969,0.00487656942965797,0.00244440185090822,0.00200331754462657,-0.00306884462326562,-0.00718106222110859,0.00653585802039114
"2184",-0.0151366880933741,-0.0211885508371822,-0.0320134021902402,-0.0298823462190841,0.00913071952890543,0.00309438126127315,-0.0189943715682334,-0.0218061013364784,-0.00324553053581345,-0.012337627793219
"2185",0.0251310061567065,0.0291119714684422,0.0234988842117627,0.0317361151622353,-0.0147538865218716,-0.00439382135340782,0.0151403995425241,0.0251773081771289,0.000279086431837161,0.00723212063576195
"2186",-0.0133717538323048,-0.00531929107056528,-0.0017007856776059,-0.00512659012253336,0.00479841831264993,0.000375125106316432,-0.0121899326465241,-0.0138147147952223,-0.0129278277416619,-0.0130548529148178
"2187",0.00544146549697566,0.00947984998174656,-0.000851783507753501,0.0103062885245802,-0.00675170118810375,-0.0022522938925178,0.00116154935889612,0.00985747288358785,0.00235560168724014,0.00859783403115144
"2188",0.00454449204390039,-0.000963172372844823,0.000852509661423362,0.00390036898757851,0.00630028474237232,0.00263440023464856,0.0163860958270159,0.0020548989709066,-0.00206799216209796,-0.00131145753062911
"2189",-0.00371042623511175,-0.0106049436443361,-0.00255530401837345,-0.00149453139674038,0.00156547283831809,0.000938064160158847,-0.000570678990139073,-0.002819571775177,0.000565156346452156,-0.0124754099800847
"2190",0.0124992396888526,0.00682081849821969,0.00768580740654823,0.00957796014661749,-0.0191644146179469,-0.00787410871697158,0.00842281290740554,0.00385592362773757,-0.00301260588389562,0.00332449124458023
"2191",0.00866666254388537,0.016453167435007,0.00847429160280089,0.0243107033624417,-0.00377354997717394,-0.000283412932517768,0.0128821391447509,0.00717038770591616,0.0133144095691329,0.0165673099142225
"2192",-0.00224797064642257,0.00285633669657437,-0.000840170505177262,-0.00231532718844873,0.0122053794686396,0.00831673587229709,0.00978363141498284,0.0010169657932102,0.0102507317165359,-0.00651901687994838
"2193",-0.0163413861776444,-0.0256349079363927,-0.0319595473540247,-0.0185669447765276,0.0153845435477455,0.00468643587458373,-0.00332185743337254,-0.00787739730665116,0.00737934665144002,-0.0150917261893305
"2194",0.0051675574073764,-0.00219280884732886,0.00608163003546935,-0.00177353624486498,-0.0162982392089778,-0.00569047679895507,0.00874839070780431,0.00438235816157717,-0.0062265360885132,0.0113257646300211
"2195",-0.0129796586075291,-0.0302731867498141,-0.0146805100975669,-0.0186556672515464,0.013904074933943,0.00497216876601203,-0.0132156768907584,-0.0148869017707549,-0.00681837286297216,-0.0059289081563676
"2196",-0.00159861963278607,-0.00377655261811738,0,-0.0159926300196256,-0.0000821767910179627,-0.00111984036302482,0.00460400177721976,-0.00338751437014706,0.00398923829678788,-0.00795224601006539
"2197",-0.0036159291247766,-0.00404334848278121,-0.00701137399287621,-0.00429326637575789,0.0068161406403342,0.00149544960547243,-0.00916560113715137,0.00967328667112466,0.0209757621421571,0.00601201054571754
"2198",-0.000259067809863511,0.00659726956566642,0.0247129973043283,-0.00215578476381428,-0.00864588121622334,-0.00261311102456796,0.00503664902082912,0.0137237309931681,-0.00615440322480598,0.00597601393501157
"2199",-0.0250973327335934,-0.0186537308669857,-0.0241169940942877,-0.0212964540426495,0.0171137981992435,0.00570766874079753,-0.018018135729193,-0.0153260351146324,-0.0126582280786489,-0.0138613336739144
"2200",0.000585291709331415,0.00436671623751761,-0.0123566673093308,0.00473042951860303,0.00283091871624763,0.00344222040231279,0.00702429380860581,0.00337254261630027,-0.00405824578598513,0.00669341801839107
"2201",0.0186582579332302,0.017902602167261,0.0214478094082964,0.0288762084866239,-0.00346815395034061,0.000185914124621211,0.0099640869302573,0.0170630626239185,-0.010372309398806,0.00731379861976911
"2202",0.00260925767100861,0.000251600737514179,0.0069991771799216,0.00549124441776305,0.0042661142477356,0.000779518335629614,0.00465104766042823,0.00152488393867567,-0.00121652628470403,-0.00660057038275963
"2203",0.014937783455649,0.019844016031096,0.0121631652025951,0.0266989228737373,0.0060580044721934,0.00482445360230166,0.00869844371757456,0.0114213764143247,0.0211748799444895,0.00664442739342297
"2204",0.0177947409184409,0.018965602722284,0.0248928333927727,0.0215722128459046,-0.0135678033274456,-0.00553959631060608,0.0179413356268319,0.0225847699224131,-0.00201854302263582,0.0132014125057576
"2205",-0.00342617701645309,0.004592798283932,-0.00837518016007721,-0.00173557233095989,0.00431361381563211,0.00204230295133478,-0.00245930951328155,-0.00318991157711679,0.0100211825876946,0.0195439748149826
"2206",0.00819068290766611,0.00962438190086234,0.0160472431428358,0.026659019508589,-0.00332305053950954,-0.00250138104346442,0.00972476783928311,0,-0.0014564354500598,-0.00191690668555067
"2207",0.00902645376664957,0.00881825817603077,0.00332488672368747,0.0107253271370606,-0.00837436197868002,-0.00260098543052967,0.00827475650928156,0.00960104644414228,-0.00510481326631207,0.00448137263945814
"2208",0.000596386625113965,0.000944887320400101,0.00248559926099445,0.00363044088866515,0.0026238479412839,0.000558717522912255,-0.00107630565391736,-0.00414525760806339,0.015851237088613,0.00446151072916767
"2209",0.0009437540670445,-0.0035403505271645,0.00165290494236503,-0.00751291005783272,0.00760546037762078,0.00335059690801964,0.00538716411708795,-0.0019589691216797,0.00396856668254975,-0.0158629878376184
"2210",-0.00630216935745709,-0.0106583224214746,-0.010726164076077,-0.0162598645934248,0.0017043269614605,0.000928139073661738,-0.00736765582583743,-0.00981335339349521,0.00494118237249452,-0.00644743147882887
"2211",-0.00479412630628517,0.00526696849443131,-0.0116763943200718,0.00769444907302907,0.00875073584925667,0.0054677445243847,-0.00647792737989994,0.00941515005518934,0.01743247794178,0.00259568152702783
"2212",0.0153547856046459,0.0126218880548916,0.0253164860228656,0.0243213156358575,-0.00489965452546004,-0.00341070514499309,0.0114099887157146,0.0130092884276907,-0.00456899226024055,-0.00258896140772769
"2213",0.00454652840033698,-0.00188162930482227,0.00493839870053447,0.000828145084889265,0.000322776044704653,-0.000832294689280699,0.00805802189454008,0.00314991169054535,-0.00706154994208186,0.000648920381757012
"2214",0.000491789576133383,-0.00376980878896793,-0.00491413076355751,-0.0102067694174532,-0.00274330697125769,-0.00046257774910663,0.0118570312882673,0.000966251688571784,-0.004178158132779,-0.0181582545830651
"2215",-0.00127820089285446,-0.00307472061663971,-0.00576119179246093,-0.000278978616932046,-0.00614944616488333,-0.00342657966907944,0.00118522373191765,-0.00120660857640242,0.0063382076326961,0.00198147886929001
"2216",-0.0062036354074162,-0.00450794364374529,0.013244973100714,-0.0144966894398717,0.00993254123302223,0.00343836148865129,-0.00355125556212599,-0.00507391033099835,-0.00887075289086969,-0.00856956398348829
"2217",0.0168936070703283,0.010247922411218,0.0122548262522428,0.0206507388475732,0.00169279507872022,0.00101847595777316,0.0109545356661847,0.0179703353385006,-0.000358014847632204,0.00332449124458023
"2218",0.0109618051968456,0.00825667680786468,0.00968541327341943,0.00582044793745595,-0.00853056787654127,-0.00564328357565314,-0.00913849430155134,0.0023851721381114,-0.0017011549520789,-0.00596420155884292
"2219",-0.00245781016918345,-0.00491346444029295,-0.000799551879113958,-0.00909354773358728,0.00665625126229319,0.00260510637959244,-0.00013151677131451,-0.00380756799983495,-0.000627802690582935,-0.00266663025528879
"2220",-0.00193234864122682,-0.00940495792276586,-0.00800006044951151,-0.0114015418706392,0.00249918442900565,0.00250540850162095,-0.0025037279650213,-0.000955601716360333,0.00224356097998735,-0.00467914912177814
"2221",0.0113745700525427,0.00735795608657774,0.00967758112823036,-0.0115330679996879,-0.00402122450920517,-0.00518376902439521,0.00383088686135813,0,-0.00805874820916908,0.0167897693851011
"2222",-0.000574215591526928,-0.00424108250748634,-0.0111821047948581,-0.00939092188732871,-0.0159092137389107,-0.00614099206389973,-0.00105261930643807,-0.00645638602564924,-0.00956849620480682,-0.00594450458779516
"2223",-0.00430968550223099,-0.000709798440361897,-0.00484658482757161,0.00172360616456313,0.00754985968357635,0.00196599308511014,-0.00724556990485681,-0.00216601793866711,-0.00382790736576821,0.00996670947658385
"2224",0.0118308732578043,0.0113662911666976,0.0073051721258568,0.0197877373155784,-0.00459559278434463,-0.00287305293282047,0.0221603043747991,0.00554743413131531,-0.00649594675674436,-0.00526308626300498
"2225",0.00289938591054129,-0.00210728399284532,-0.000805884833434911,0.0132170783875116,-0.00820009021207146,-0.00262784991384779,-0.0098664160160068,-0.0040775181990258,-0.0148263473552389,0.0178571708144006
"2226",-0.00303330471614138,-0.00680418724551035,-0.00483850437150413,-0.00804887178436287,0.00115739953802052,-0.00103487902812638,-0.00432654798437138,-0.0144507643142596,-0.00944103544285746,-0.0168941229624917
"2227",-0.000998236630679439,-0.00307108840684855,0.00729333156653467,0.00167881909011136,-0.00264262937716409,-0.000659652391510668,0.00289708962893087,0.00171032848640085,-0.00311410773696219,-0.0079312219733344
"2228",-0.000523392020839841,-0.00545037266904314,-0.00241369834258931,-0.0139664594098798,-0.0146557877837228,-0.00678669441662882,-0.028623930842881,-0.0124419409016485,-0.0145778210391692,-0.0059960575746596
"2229",-0.00933154702885208,-0.0104836577402363,-0.00403203560834886,-0.0249291749032826,-0.00563029474123555,-0.00170847283434228,-0.013517259927331,-0.0249505713333704,0.00288188286036273,-0.00871308670317672
"2230",0.00230670517186815,-0.0043343173892253,0.0105261394232989,-0.004357888709701,0.00295784069025684,0.00190135942722347,0.00918062366496919,0,-0.00210729881020499,-0.00202843934733932
"2231",-0.00393152473431391,0.00507871638952495,0.00400662650452199,0.00204265297208273,-0.00210616325013147,-0.000474161771560566,0.0012219088829768,0.00810765832959381,-0.00335955077750061,-0.0101626021929274
"2232",-0.0139598632238876,-0.0153994945446108,-0.00957719451457539,-0.00960999163178755,0.00481265785678286,0.000569545398735105,-0.0071873986010097,-0.00804245286959537,0.000192584027880471,-0.0143737315317003
"2233",-0.0112282477266686,-0.00855328664844279,-0.00483467108543911,-0.0138193796315157,0.00571417632290405,0.00379504754122295,-0.0105176475130944,-0.00481372632248445,-0.00279248922084718,-0.00763885608064085
"2234",0.0152068078206464,0.0125708747767903,0.00971667103256335,0.01937984613455,-0.000918958877485609,0.00132331696886956,0.011733831536185,0.0132381389797933,0.00144844537366651,0.00489846340708389
"2235",-0.000729291308129598,0.00316462163794284,0.00240553972466917,-0.0029246492519408,0.00167257900556139,-0.000283320464031789,0.000546020005109726,0.0047735132771074,-0.0132099413095164,-0.0153202689780357
"2236",0.0158659865649613,0.0101916586239095,0.00480012362449256,0.0108533867203449,0.00208742759595681,-0.000472061669513857,0.0106364933772893,0.0072522196254845,0.000879460655831998,0.00424322340568328
"2237",-0.000862347849295508,0.00576512480788804,0,0.00899620120890865,0.00666527830330366,0.00217268344016897,0.00283380431209213,0.00571004491167848,0.0110319047154153,0
"2238",0.00364409123437448,-0.00740386712927976,0.00477695343181117,0.0100660700826243,-0.00306268658133935,-0.00131985489263076,0.0102260047699365,0.00444341467728049,-0.00453845122708474,-0.00140843151233594
"2239",-0.00114685288744176,-0.00697792418724918,-0.00475424263613489,-0.00939642928235052,0.00307209544684106,0.00132159921181652,0.00173168642931132,-0.0105676759174597,-0.00805115949369128,0.0077574441065984
"2240",0.00133957455936162,-0.00169631757214028,0.00477695343181117,0.0051739210048598,-0.0000823293833634997,0.000942697326987263,-0.0049194925668935,-0.000745382379443327,0.00664971627909816,0.0160951672652541
"2241",-0.000143179038258556,0.00582529584004643,-0.00633910554705042,-0.00772078883703498,0.00231725732340449,0.000564748706982421,0.00334008289299437,0.000248745283969898,-0.00466293948585716,-0.00137739162486072
"2242",0.00114655967574384,0.00482640541036283,-0.00478474669878037,-0.0219020828554293,-0.000990840853773545,0.00103561127936702,0.00799041668879585,-0.00472164771042072,-0.0118094769842814,-0.0151724188841127
"2243",-0.00415163649706196,0,-0.00801270616668015,0.00147316231053773,0.00396776865330617,0.000376055593562352,-0.00634135465612484,0.000499195182228629,0.00661726419753084,-0.00630257884926444
"2244",0.00953554299507475,0.00696440725922698,0.0153471952151034,0.00764936803724137,0.013507601548078,0.00531820936241623,0.0123652214565266,0.0187173813067565,0.00353219198454058,0.0112756100009341
"2245",-0.0102049914280966,-0.0114476433189787,-0.00795518410948981,-0.0119710484853386,0.000325564430034175,-0.00280882396720539,-0.0189127037436239,-0.0142086974032248,-0.015545532025279,-0.0209059238447552
"2246",-0.0140028064503899,-0.00506626848801828,-0.00962316589526724,-0.00561453392174394,-0.0271832195066187,-0.0105165939467207,-0.0147256623017438,-0.00670969425222101,0.0106266757249642,0.0113878176129558
"2247",0.0195030376400305,0.00994165317987905,0.00566789232277776,0.00683502885658216,0.00878441713632183,0.003700606239881,0.0167122079295063,0.0085062639723239,0.0222090699251363,-0.0014074403706511
"2248",-0.00605848102299111,-0.00672264350000695,-0.00241548808374525,-0.0165288994772951,0.00970296243426061,0.00321517440296426,-0.00267302732591579,-0.00868267037304604,-0.0129782641697249,-0.0288936282311872
"2249",-0.00671955878386998,-0.0157117712358962,-0.0129135832525931,-0.0111043374623248,0.000492780131175818,0.000565320476173525,-0.00241148502230382,-0.0102601105820607,0.00165577094878278,-0.00507975678233286
"2250",-0.00777978179927297,-0.00221038109972982,-0.0114471903126192,-0.00819424837976168,-0.00106712447099966,0.00150685877109069,-0.0061786691355209,-0.002781426450985,-0.00194473947665263,0.000729459707354385
"2251",0.00258110091303143,-0.00319958660731645,0.00909834917361141,-0.00673205676055311,0.00131469474770962,-0.00216303397266382,-0.0056766197713215,-0.00329616780794695,-0.000876812167544982,-0.00364433985582713
"2252",-0.0193811845507025,-0.0170368380458027,-0.0155737417885333,-0.0280345681059826,0.015758626798964,0.00801142445112912,-0.00462129154495139,-0.0167896046901449,0.00546073119081236,-0.0102415653600367
"2253",0.00505246000368853,-0.00150699100638307,0.00915902297208815,0.0161649610811414,-0.0129281942845739,-0.00738670723284807,0.00314056352855641,0.0049160265520547,-0.0128018619648738,-0.00665179463204035
"2254",0.010497805170921,0.00905629000302288,-0.00412552222206553,0.0152837602038263,-0.00589385392975816,-0.00254338975263191,0.0110263482114805,0.00334698391447064,-0.00265255916443108,-0.00223211243083221
"2255",0.014632111250255,0.0184492165142276,0.0248551331748899,0.0196621758145552,-0.00214096360232463,-0.00264447551561631,0.0196583403227313,0.0207850725964656,0.0121158691523602,-0.00447421180545382
"2256",-0.015238160752032,-0.0141981294137512,-0.00970096171466772,-0.0129559054698459,0.0113056007837971,0.00416633678869016,-0.00488596822764276,-0.0145802350129201,-0.0218978102189781,-0.0104869787599111
"2257",-0.0178150946784295,-0.0124162027406515,-0.012244845477186,-0.00335751650185212,0.00554865082597789,0.00358371992362394,-0.0127388387105744,-0.00282349276230665,0.015323393034826,0.00454210752137274
"2258",0.00824906317787488,0.00475434154865395,0.0031634748368714,0.00780741063940105,-0.000243749692887429,0.000469665038589362,0.0051073508655235,0.00360395559204485,0.0108780967181683,-0.00452157006397669
"2259",0.0090744162095171,0.00729930699009995,0.00746884969450479,0.00802459373312892,-0.00722383728439657,-0.0028176554506687,0.00414560447063361,0.00487304655228082,-0.00523510411565486,-0.0045420296094798
"2260",0.0123834961479519,0.019490235988723,0.0107085205413415,0.0140844835697862,-0.00752191974616856,-0.00226035946824243,0.0113198627990501,0.00995406085308681,-0.00292372085641046,0.0182510150888562
"2261",-0.00165066240365563,0.00147066260699957,-0.0122250286243372,-0.00362312412319232,0.00572924903505045,0.00183428929516904,0.000266598366961412,0.00151622355868097,0.0072329685706769,0
"2262",-0.00228492247560164,-0.00416049135006047,0.000825158700619166,-0.00696965140533956,0.00295457889984196,0.000188455547719846,0.00293359602261734,-0.00656054408575324,-0.00756919919740318,-0.0141898071176862
"2263",0.0106717693710769,0.00884706701167559,0.0148394266702847,0.000915353433573518,-0.0166130012162087,-0.00528333918880874,0.0102365233880408,0.0104137844802918,-0.000684462716861178,0.0166667524346811
"2264",-0.00708776702787939,-0.00803867159684757,-0.00568662722067526,-0.01554870793412,-0.000998851775883991,0.000379464380007688,-0.00447438067835149,-0.00703846893517734,-0.00763208437276164,-0.00968705542198245
"2265",-0.0100033693351818,-0.0149805030807205,-0.00980398495091306,-0.00309707382270319,0.0044986692270943,0.00113763969038105,-0.00753461325949834,-0.00962059123286918,0.000394409394486317,0.00526712378627625
"2266",-0.0139795430994832,-0.0149589902243605,-0.0156765395781253,-0.0273376711147233,0.00721488377095181,0.00426188396039495,-0.00972295142514845,-0.00894701082068339,0.0140942244637712,-0.00748492787745059
"2267",0.0016913860447878,-0.00632723723389206,0.0125734148845289,0.00223586895484851,-0.00403469429767289,-0.000282961103952095,0.0164091477995516,0.00154805615773457,0.00281855382270924,-0.0098039421145949
"2268",-0.0126141759479956,-0.0168112375105918,-0.0173842065402128,-0.0191203655555258,0.0134757689769742,0.00603680827885777,-0.00330864514418505,-0.0100439872193487,0.0144407637138981,-0.0159939228439159
"2269",-0.0239914291558162,-0.0181345931099194,-0.0151642189563559,-0.0308644499274063,0.00179468741273348,0.00215680741487412,-0.02230469672046,-0.0228927783025503,0.0141397155658682,-0.00464405853976857
"2270",-0.0109765890671502,-0.0100264983517603,-0.0213858261838878,-0.0107274645696325,0.00447807410148537,0.00252663556421084,-0.0118141172616196,-0.0135782234734825,-0.0044277154135145,-0.00466564641415823
"2271",0.000990126800631597,0.00346488724518745,0.00699308402258869,-0.000338812004883726,-0.0109431711141263,-0.00317351733105864,0.00398509792307244,0.00377858186543945,-0.00889479560938689,-0.027343700059397
"2272",0.00806820393644347,0.00796825628412523,-0.00520836678174919,0.00203386225901858,0.0144246931480043,0.00449372589719665,-0.00698077284392129,0.00430224010495972,-0.00506013948940498,-0.00642569783124736
"2273",-0.0249406536055898,-0.0171277113193101,-0.00872602829326719,-0.0104870595153169,0.00985709984792726,0.00391523194872856,-0.0151618869783308,-0.0109771020153471,0.00489398334990865,-0.00565877484512667
"2274",0.016416701311222,0.0128684808198591,0.0123240553375761,0.0129915005882701,-0.009360594301425,-0.00204302724387173,-0.00139949923667537,0.00893345500086062,-0.0162338042758421,0.00243899091980437
"2275",-0.021466010294429,-0.0367921261965688,-0.0278261071200259,-0.0394870525431716,0.0155870359394059,0.00465162867016389,-0.0113524086242407,-0.0300511378591172,0.0102893130544353,-0.0210869089061161
"2276",0.00133107130069154,0.00906861715744323,0.00805012877510602,0.0147574873455842,-0.00310138482649314,-0.00129672223683364,0.00297729427907512,0.00553250482299705,-0.000960789758632008,-0.00828489181420122
"2277",-0.0128150304926715,-0.0206971504519684,-0.0381545183317613,-0.0218143643579174,0.010529625864232,0.00491486328876922,-0.0265730945308066,-0.0220080403632341,0.0133679549903456,-0.0075187801837816
"2278",0.00560205041996076,0.0108454686123984,-0.00369002749083225,0.00389398523744244,-0.00678879997497051,-0.00249120134932423,0.00667974204337551,0.00450063644800669,0.0011387965890064,0.0134680023834841
"2279",0.020515116335994,0.0264097193468225,0.0453703420716749,0.0342029076331489,-0.00381494514648539,-0.00221965707911553,0.0276935654041712,0.0229626059690105,-0.00464497117537155,0.0299002652026497
"2280",-0.0151163930900197,-0.0134012033175865,-0.0212578884163688,-0.0170473292392546,0.00542545421810869,0.00333692280878206,-0.00982459415240244,-0.00848612171427643,0.0102857333333333,-0.021774146157322
"2281",0.0136429952627484,0.0214613191670312,0.0135748611593092,0.0145681300232499,0.000475691190758631,0.00073907217515301,0.0214032129389619,0.0168415983012167,0.0114064760292898,0.0197856396611851
"2282",-0.0108832462620551,-0.00851055162185044,0.000892721751707848,-0.00341872999818127,-0.000237599230065166,0.00073874862207024,-0.0155424513487386,-0.00705945242821859,0.00372822253958227,0.0121261125018888
"2283",0.00520920521908996,0.00214624720592549,0.00178409276779568,0.0157804183860617,0.00142796937644452,0.00129177496575816,-0.00662555763169703,0.00710964261201985,-0.0106788093475939,0.0111821204449172
"2284",0.0243775216350479,0.0160598753691636,0.0240429859899869,0.0324214267021363,0.00847672130236798,0.00534369786586431,0.0217114952019908,0.0285094333786804,0.00384828229915257,0.00947862482423667
"2285",-0.000361501760742566,-0.00158069096615909,-0.00608697566067506,-0.00948641349748558,-0.0030618707454908,-0.00230352764483899,0.000138857671614812,0.00712769027501547,0.0102852363801376,-0.0187792482003014
"2286",-0.0180222008895534,-0.0274405362492751,-0.0104986599097435,-0.0323645841549108,0.0185524623790312,0.00708344501037761,-0.0105540183130968,-0.0212320839764264,0.000370134186854276,-0.0175439474833902
"2287",0.00599487034842894,0.0151926709440655,-0.0123784410226562,0.0283276844117439,-0.0082934433243097,-0.00109608081089096,0.00491209635717538,0.0182111300801779,0.010731834979437,0.0251624127265246
"2288",0.00156831935373591,0.00133617451074297,-0.00268606157392337,0.0076336114261808,0.00484575157378653,0.00237792061305098,0.00111751687181827,0.00236705559139549,0.0120823798627001,-0.00158359108553852
"2289",-0.0190499673041427,-0.0152123392467303,-0.0170555542338099,-0.0115285355705117,0.00116669586703821,0.00127766884361979,-0.0224610752185594,-0.0170557826092083,0.0158270778692231,-0.00634416643820135
"2290",-0.0134612385958759,-0.0235772618046641,-0.00182643002313465,-0.0136620319768538,0.0215195927682421,0.00747143504121195,-0.0293989279654422,-0.0149489710512868,0.01344375,-0.00478852442938482
"2291",0.0000538343352312065,-0.00888149109875036,-0.0192131139997107,-0.0138513059764714,0.00106450210648679,0.000180648514132908,-0.01617406382124,-0.00406555033788447,-0.00219625753850028,-0.0256615684840983
"2292",-0.000862639426941647,0.00420044340764725,-0.0177239739338021,0.00411096191310545,0.00881285507681095,0.00298363018347958,0.00523085257225731,0.000272215020091338,0.00774781638056332,0.0016460680853132
"2293",-0.0130081961606465,-0.0142218466941039,-0.0199430604897948,-0.0167178377785114,0.00700327422297553,0.00459818091062436,-0.014719110247802,-0.00843295387347698,0.0401887038283129,0.0123253916243458
"2294",0.0206169737245514,0.0195191558800756,0.00872110588135011,0.0173491150670153,-0.0166018544977853,-0.00762812589857009,0.0129770666878057,0.0150889202895204,-0.00587936344497497,0.0146104412805887
"2295",0.016878297924575,0.0160929591834036,0.0365032406167609,0.0221692027042228,-0.0105701794218857,-0.00298458214901298,0.019216638059526,0.0202705364565243,-0.0303312265095367,-0.0112000939303752
"2296",0.0163347844637616,0.0207537993959095,0.00834099801588506,0.0196861626671199,-0.00614885514925323,-0.00244893717278349,0.00906159133478956,0.0127150789808066,0.00618633805488367,0.0210357295389787
"2297",-0.00409589150193357,-0.00588542977610873,0,-0.00588991210112844,0.0122960769939933,0.00463732274474116,0.00955966748946624,-0.00392328412923793,0.0243331999220679,-0.00554667519181595
"2298",-0.000468424890686991,-0.00188370220003686,-0.00459544002389967,-0.00460833486443579,0.000840353677504124,0,0.0021520583394492,0.00787792497527962,-0.00600218948345443,-0.00876506550734024
"2299",0.0144789704480619,0.00727972590345538,0.0166205056158337,0.0248016247997735,-0.000534329261787092,-0.000995196548846056,0.0115964016995229,0.0104220962406121,-0.0177751655421812,0.015273351601643
"2300",-0.0126296014072507,-0.0173985338315223,-0.0163487806157969,-0.0212972082919769,0.00404770964467294,0.00199275207731686,-0.00240591985107785,-0.0167615175265198,0.0149796781536007,-0.0134600760332335
"2301",0.00457568325137214,-0.00435836214464036,0.0101569575820042,-0.00230792934894919,-0.00197760289538595,0,0.000425412069969378,0.00550778703565435,0.00332707726218162,0.0128411642829631
"2302",0.0121118801312277,0.0139533609574434,0.0118828560876694,0.00330476850707262,0.00358180166810551,0.00298381566731987,0.0181512296586321,0.00834604471119005,0.00263580475609393,-0.000792463724620274
"2303",-0.00230139272547447,-0.00296810871014963,-0.000903230004450806,-0.0098815026080461,-0.00964463136177207,-0.00486778022084455,-0.00306445641207753,-0.00646618219153616,-0.00686903844757536,-0.00158593958574915
"2304",-0.00784253618828457,-0.00460087382295593,-0.0153706293216243,0.00864941127605845,0.00437109012919112,0.00163083402247777,-0.00167641906937055,-0.00104159502418,0.0130646228924549,0.012708406021543
"2305",0.0235071992574138,0.0274607034146381,0.024793261125178,0.0356199676570121,-0.0176089802145424,-0.0078165268071968,0.0260288384190448,0.0242377715128743,-0.00733312548325293,0.00078430302575816
"2306",0.00449217153157644,0.00238168761307,0.0143371731000326,0.0133758065883236,0.00412716427535953,-0.00173440209676468,0.0076374650076303,0.00585221118897605,0.00772695103320764,0.00548589929572096
"2307",0.0039196788994369,0.00844761015197304,0.00706683107548911,0.0113136130004912,0.00364439540946382,0.00118880469229699,0.00500830302612654,0.00455357534176559,0.0172733653522075,0.00545596840250417
"2308",0.00325360356921922,0.00523577662161268,0.0105264801901495,0.0198881795809476,-0.00641272454184449,-0.0033795295416319,0.00269351082054237,0.00302232226114718,-0.00157377615570831,0.0193798199127144
"2309",0.000798332914656141,0,-0.0104168276601408,-0.00152337782514911,-0.000310911626960619,-0.00201603079209933,0.00188035429789801,-0.0057750335812744,0.00497758416311944,0.0182510150888562
"2310",-0.0109178979322492,-0.010677187717115,-0.00964903975172937,-0.0170889815127012,0.011045556907509,0.00578502140258541,-0.0103228581606762,-0.00303008378833425,-0.00462272580999457,-0.0134429144816003
"2311",0.00493963849592194,0.00552770198139863,-0.00088589337162992,0.00620939497661621,-0.00607816619817303,-0.00392582637698347,0.00406383278422662,0.000253458527296191,-0.00829324915751783,0.0151400727276354
"2312",0.000802454282426091,-0.000523556621304988,-0.0044325775337094,0.00154271767135583,-0.00410241760237162,-0.00357443369445454,-0.0025634295171445,0.00177252192453037,0.0160561796946617,-0.00149140393515124
"2313",0.0161370784387498,0.0267154649202028,0.0267143350324748,0.0209488409694392,-0.0101040660092713,-0.00285157546827075,0.0236711373088649,0.0245199563898735,-0.0172016131687243,0.00373407885778065
"2314",-0.00128233235444641,-0.00280607417018952,0.0043363964136367,-0.00603520857880757,0.00314071002350924,0.000737925404911355,-0.00132152843519129,-0.00197399611206794,-0.0128967502588812,-0.00892852630190855
"2315",-0.00162963804919869,-0.00946524252510295,-0.0129532070304652,-0.0142680935625762,0.000939085729732447,-0.000184320172135322,-0.000264608131771649,-0.00296703040725099,0.000763519111813382,-0.00825829985097226
"2316",0.00578720257932974,0.0103304478234514,0.00174965810467675,0.0200183722144136,0.00297160399705931,0.00525524524031784,0.0127052933598901,0.0126459872634757,0.0222956682120692,0.0174110485764289
"2317",0.00634402364172182,0.00741312572683417,0.00349334630401676,0.02204102949609,0.00413203307645138,0.00110054249829883,0.0139831814762061,0.0173847378339598,-0.00381457015721265,0.0111607918898995
"2318",0.00392977517945003,-0.000253624432997812,-0.003481185318152,0.00531758182322584,0.00209672546640483,0.00174089824403389,-0.00386656109547312,-0.00166686354281786,-0.00274697417997938,-0.000735900819623936
"2319",0.00141902746091227,-0.00482250557780162,0.00436695506177465,0.00205709177165581,-0.00767067670739829,-0.00283529492009915,-0.00646930806706092,-0.00121014972341293,-0.00701171935696865,0.00294554370651778
"2320",-0.000537775599956714,-0.00535571107366661,0.00608669287982333,-0.00234594501236751,-0.000234617036095175,-0.00210939480500494,0.000260966352427783,-0.000727033370522268,0.00294215705230449,0.00734219461659547
"2321",-0.00659921680745479,-0.0082051310436182,-0.0129644738446856,-0.0170488380547478,0.0113247589231027,0.00459542407795732,-0.00704847350154114,-0.0106692756297103,-0.0226300984432167,-0.0211371111512028
"2322",-0.000442983980164957,-0.00723868529252636,-0.0061295937900655,-0.00239234608697625,0.000386048062876121,-0.00100635023801476,0.000796126240879769,-0.00661732237186363,-0.00240115768457971,-0.0059567318472874
"2323",0.00059068948816754,0.00416660748600717,0.014978091394114,0.00329724776507434,0.0013125290077991,0.00146534302899171,0.00768942147418072,0.00320684056697806,0.00232094898442448,0.00299621356440394
"2324",0.00925024111498907,0.0121886521936154,0.010416568894374,0.0137436285616732,0.010485177687771,0.00676732378821288,0.0198654109325742,0.0150029334069515,0.0185249059781287,-0.00224052417919829
"2325",0.00438770979284175,0.0107608208285501,-0.00343634763129042,0.0103155107381268,-0.010529361236093,-0.00136254630064625,-0.00154763618808762,0.00823841437891026,-0.0139778037390064,-0.00374246393872524
"2326",-0.00242688853295159,-0.00861850495245042,-0.0163793029133185,-0.000875227434378179,0.00709407726203382,0.00363806363253794,0.00594286626209151,-0.00360502063765245,0.00461145182940137,-0.00150268636214512
"2327",0.00681172238402272,-0.00869322380319359,-0.0245400034866394,-0.00291964529535038,0.00260851699601572,-0.000290544259282099,0.000642455970634614,-0.0089242357093765,-0.00603535367252084,-0.0173061642997535
"2328",-0.0032380207540551,0.00128964805180365,0,-0.0120059133117398,0.000612160815353535,0.00118077491892832,-0.0014122145020532,-0.00292023249986961,-0.00667064055417776,-0.0137825107354482
"2329",-0.00998767101377496,-0.0190625625673442,-0.0215631916332455,-0.0195613986021722,0.010936376455901,0.00399003114164143,-0.00565534803833723,-0.00610231064999578,0.0130004474730874,-0.00232932034986943
"2330",0.0109211846843096,0.0152312623173503,0.0165287329148496,0.0120919077669168,-0.00726254628475453,-0.00216791649309167,0.00245610053882395,0.00982320430558037,-0.00611934366413924,0.0108950335716682
"2331",-0.0119659376325956,-0.0168131585093853,-0.00541989411576849,-0.0200119461132946,0.0123450363329076,0.00515996713727152,-0.00541587518732789,-0.00851177171497419,0.0142808189792916,-0.00307932878634831
"2332",0.00269664098012212,0.0176268485483158,0.0290645098120104,0.0173727823712351,-0.00632292174947358,-0.00153110132536016,0.00570445746820836,0.012999832746007,-0.00151758703720095,0.0239382940858939
"2333",-0.00234698018104074,0.00180967874447102,-0.00617828350950544,0.0128819247633378,-0.00128808337277397,-0.000180376885494105,-0.00128912357269784,0.00411618400205316,0.0135100819049228,0.00754137452184356
"2334",0.00931272497538327,0.0113547023960574,0.0230905737058651,0.015380142652653,-0.00690241478249454,-0.00396938087584986,0.00684159820013686,0.00795775207867666,0.000166658336804515,0.02170659899314
"2335",0.0101009470526172,0.0137791973103003,0.0277778228657524,0.0177688086619752,0.0035133529186484,0.000724523446614889,-0.00230796794697496,0.00885151955048458,-0.0106622737860324,0.00512828594201653
"2336",0.0000481495929676168,0.00125860185977356,0.00422292742820662,-0.00486540714594275,-0.00479482462663239,-0.00235308267881984,-0.00642495646819508,-0.00545398582834633,-0.0139765600903401,-0.0080175326796712
"2337",-0.00110585966924737,-0.001759666040134,-0.00925145907757685,-0.00575227984597371,0.00856568110672562,0.00299400277301443,0.00659595905145904,-0.00238433215927791,0.00691654848504375,-0.00367379462428574
"2338",0.00702675300293687,0.00906551902705344,0.00763994435286319,0.00462832590334306,-0.00432265149490763,-0.000995169638337234,0.00424007602341825,0.00693119625407879,-0.0015264586419006,0.00442479420991582
"2339",0.00315425391195712,0.0197156803248213,0.0151642874479381,0.0152604801798368,-0.00312198626907867,-0.00162951578349457,0.00102338420168246,0.00593397885701119,0.0156276883918411,0.0212922283683834
"2340",0.000952761031621563,-0.00244733628174842,0.00580912530860633,-0.00453756585353715,-0.0110004243720676,-0.00507857623684216,-0.0140592580599449,0.00259542948833702,-0.00510119576683066,0.0194104523215852
"2341",-0.00537817669389795,-0.00711485345524243,0,-0.00997146881261624,-0.00594839786786427,-0.00164073527963371,-0.0169818868901296,-0.0112967384234534,0.00378244091970714,-0.0042313265506686
"2342",0,-0.00222382576509561,0.00742580223675593,-0.00604344074858987,-0.00256417900902373,-0.00109583002701397,0.0106814718300789,-0.000714038881167167,-0.0128119161415494,-0.00424916097384553
"2343",-0.00172293750068353,-0.0042101746722023,-0.00655198975595184,-0.00636936796244547,-0.00412908524561684,-0.00109649447088067,0.00626323954289232,0.00905204229746825,0.00288407840261318,-0.000711300967053075
"2344",0.00148618754233598,0.00547121006186146,-0.00412198973459177,0.0107808783212238,-0.0045372423108182,-0.00210443223404233,0.00363084245624079,0.00779033690939346,0.00397525152731326,0.0128112856578488
"2345",0.00205819951897435,0.00469953415328805,-0.000827868499405082,0.006053734773243,0.00998042782396769,0.00550121378040025,-0.00025876523093038,-0.00163990113413781,0.00286439771350633,0.00913564938547906
"2346",-0.00907586651739134,-0.00516980371943887,-0.0455674627933527,-0.0103153526101952,0.00412387530742375,0.00346572233906972,-0.00232588271698686,-0.0063351757662331,0.0189012095186389,0.00557102644813079
"2347",-0.00539883876834479,-0.00247473170326951,-0.00868067403401029,-0.00434261785837609,0.00255749154238516,-0.000363712357860035,-0.00829037628996998,0.00023645442817255,0.0194575066414584,0.00969530142169384
"2348",0.00794846569982277,0.0074422432768031,0.01838863898927,-0.00261712240503542,-0.0100683027179047,-0.00290429993194941,0.0133228736687532,0.00873419075114601,-0.00331584305190713,-0.0137173754198485
"2349",-0.00870316135919014,-0.0201917099844675,-0.00945803068932261,-0.0282798567847307,0.0125956886919771,0.00593510151488608,-0.00219133533780791,-0.0109991242697192,-0.00227198153638397,-0.015299103572847
"2350",-0.00557836353974706,-0.0130686913287327,-0.00868067403401029,-0.0162016989659498,0.00548549139882204,0.00181538688926586,0.0134350864029269,-0.00567864353746528,-0.00609954461694495,0.000706277775116781
"2351",-0.000194755307658112,-0.00483844072251505,0.00525387990396697,-0.000304852713861603,0.00668498995489597,0.00271781564953177,0.00382400377016912,-0.000238373929529856,-0.00114556092910212,-0.00988003858289233
"2352",0.0036588979865404,0.00307057404782429,0.00522660976519052,0.00152527057278617,-0.00427407377619815,-0.00234904151138182,0.00977801024250602,0.00166622650928949,0.0090931432784469,0.00641481120450282
"2353",0.000826320657348445,-0.00127538440723407,-0.000866513683326353,-0.012793119041549,0.0031428885264877,0.0019016556486986,0.00804816359627458,0.000713007525933396,-0.0205390323104401,-0.0219545936385844
"2354",0.0124339590252649,0.0102169845879145,0.0251517949103408,0.0191296374325576,0.0000758811810441795,-0.000180746169438195,0.00187127315598601,0.0121110849005437,0.00273519266083389,0.0246197266652655
"2355",-0.00935480175892678,-0.00581544224059172,-0.0186125412845435,-0.00242187473989186,0.00565464693740325,0.00153727428329109,-0.0178061212526041,-0.0114968047683649,0.0094230448977588,0.0233216012391908
"2356",0.000290513187308328,-0.00279753962290463,0.00775858888924108,-0.00273136282534991,-0.00455890049683205,-0.00270845346747206,0.00494423113560538,-0.00617157423183801,-0.00786111182784688,0.0013812676985363
"2357",-0.00871432852347898,-0.0102013516370694,-0.0136868768298618,-0.0179549568890988,0.00969392802101132,0.00380222138374209,-0.0080736663461134,-0.0100306934358491,0.00453941054673446,-0.00137936242976755
"2358",0.00986543646888927,0.0123679203187281,0.0138768069777582,0.0120855200876415,-0.00861793375531583,-0.00360706196799354,0.00788500801807346,0.0123039241622547,0.000739495528218725,0.0110497861959944
"2359",-0.00933348064799377,-0.00865362966793759,-0.00684353114319236,-0.00459279447759975,0.00167745864130153,-0.00135776652079234,-0.0151419951587891,-0.00166830573304921,0.00344825935677506,0.00751355819875688
"2360",0.000292607080950136,0.00333758949668539,0.000861312630645594,-0.00984320109556447,-0.0142354725166083,-0.00806592434462694,-0.0139651033495601,-0.00405827147507887,-0.0173457943270676,-0.00745752564579838
"2361",-0.00346503981876078,-0.00614129500322658,-0.00688459459868529,-0.00931960335584814,0.00432443216882317,0.00100485456564758,-0.0107848660026884,-0.0105466161037607,-0.001915029174272,-0.00273227328300718
"2362",0.00631756497845215,0.00823893228829831,0.00693232081713946,0.0100344317712768,0.000769025023747094,0.000639154013448051,0.0080125679113412,0.00436044240428179,-0.00133481268036673,0.00410953283883031
"2363",-0.00136262460506642,-0.00306418401582775,-0.00430299697841485,-0.00186260467796917,0.00222819580043976,0.000638448060862329,0.000912239928324787,-0.00024092696299749,-0.0028401637527371,-0.00545702180239194
"2364",0.012962225797283,0.0197232237531035,0.00777880141933829,0.0102642025790123,-0.0044459045442653,-0.0016409821044947,0.0119774910419281,0.0125451314959486,-0.0173410400266136,0
"2365",0.00678305453878125,0.0113035579111105,0.00686113952862422,0.0120074507281869,-0.00377392341943239,-0.000456676929605271,0.0015435759446758,0.00309693910580511,-0.00272804767106449,0.0116597902841575
"2366",0.000286811243185081,0.00372595719184843,-0.000851775051887382,0.00669310606391882,0.00517905690908282,0.00310621573575554,0.000642417548623708,0,-0.00341939639033861,-0.000677887099525876
"2367",0.00429934386799546,-0.00247473170326951,-0.00255754977942735,-0.000302256676409929,-0.00146101352374062,-0.00191257112650656,0.00436453112317259,-0.00118732307175851,-0.00823467990676474,0.00407050060119052
"2368",-0.00190260696639588,-0.00843463163332681,0.00769234599910895,0.00120919077669179,0.00238727058363941,0.00118636426530516,0.000127933364223676,-0.00784764488632861,0.00380552662673783,-0.00608106773660633
"2369",0.00204925405389544,-0.00125092975867824,-0.000848139749268562,-0.000603865200115461,0.00405728510570857,-0.000337655960163108,0.00063913347197464,0.00143806735560914,-0.00103391351083759,0.0101970756409457
"2370",0.0030435375930451,0.00300610675838153,-0.0084889190785421,0.00815702209646374,0.00720725012913537,0.00310406652559769,0.00536366757552731,-0.000957271842675134,-0.00232882521426903,0.00201895364593252
"2371",-0.00298697318408958,0.00549432445085229,0.00428070608703734,0.0152832513967347,0.0142355205726306,0.0092835118657919,0.00304898592747183,0.0162911698911015,0.0277513534667821,0.00671589392978178
"2372",0.00508851555759349,0.00322918951860696,0.0102302453237364,0.0106257134731735,-0.00743068971593008,-0.00261532933505981,-0.00620575505359289,0.00660073605977596,0.000336482175382402,0.0120079785873621
"2373",0.00156114307690669,0.00693233308767272,0.00675096856746427,0.0090536969981867,0.00242052645892699,0.00144656717631686,0.00611706862963168,0.00491793489216885,-0.00084088464246368,0.00988800541244195
"2374",0.00325983323358536,0.0022131160014347,0.00586755726765342,0.00723597655590535,0.00535583189440514,0.0011739218850304,0.00531961320002794,0.004660744069795,0.0148123379902374,0.0169711811449773
"2375",-0.0013656393602155,-0.014475128282106,-0.0116668629899177,-0.0114941340004283,0.00645287050916199,0.00153314098238799,0.00151200814737629,-0.00347915851615022,0.00555646034903878,-0.00192551936769392
"2376",-0.00947739375949597,-0.0343540190652999,-0.0177065240352851,-0.0252907301529485,0.00484608826739019,0.00351149832137776,-0.00490615575883713,-0.0188549853331591,0.00404122061855672,-0.0122186152959649
"2377",-0.00771175919943301,-0.0152100321942406,-0.0180256034163011,-0.0140172908974887,0.00445176848111184,0.00197398778642199,-0.000758703561325347,-0.00972688991122073,0.00739281267279135,0
"2378",-0.00196690655126452,-0.0185865005232561,-0.00437067751411779,-0.00332740356112249,-0.000738289301650541,-0.000268438490402478,-0.00544021015999496,-0.012937571151816,0.00105999674706458,-0.00651046168649383
"2379",-0.00139406281110988,0.00533481187179485,0.0096577726066287,0.0106223148981766,0.00384354622850847,0.00304546796806404,0.00915909691002437,0.00339816192394604,0.00741225887624641,-0.00524239253493219
"2380",0.00298420453276971,0.00716383802266374,-0.00434796768229606,-0.00360373931735836,0.00485983118755406,0.00107149908375259,0.00504212264945902,-0.00072554770492872,-0.0105110203751617,-0.0171278363614298
"2381",-0.00372397386827461,0.0150153996148712,-0.00174660214807265,0.0027125297017716,-0.00622891105686074,-0.00338952939184056,-0.00150507770033226,0.00383304244146876,0.012828893924552,0.0234584695446547
"2382",0.00644010894454117,0.0254348880003443,0.0227470727617216,0.0177335565045331,-0.0106924756027911,-0.00429665074235996,0.00188454171476149,0.0248051179501381,-0.0059701332626898,0.00916831322138223
"2383",0.00283857844629143,0.0102058185170957,0.00684353114319225,0.00767891309484781,-0.00462158118135669,-0.00224756113924574,0.00411156141982438,0.00783102261061552,-0.0192354761726765,-0.00778717815876662
"2384",-0.00163116655270823,0.00205139913026997,-0.00924829554833118,0.00254006713197352,0.00164767853347603,0.0019822473094917,-0.000503969634002233,-0.00306120404121468,0.000496573998562511,-0.0058862543246091
"2385",0.0130224505973831,0.0307061839217035,0.022471869900327,0.0241602949458593,-0.0114382221965124,-0.00476602081450972,0.00668067407524875,0.0174776974424009,-0.00653433405236836,0.00789483252926959
"2386",-0.0359089993489581,-0.109483659624432,-0.0414200161314434,-0.0607018625910941,0.0268469742490647,0.0138235097741992,-0.0121460357298108,-0.0733519494909414,0.0490383727496597,-0.0202349783501855
"2387",-0.0179100389828449,-0.0231393235723737,-0.00529110490131413,-0.0128638213021902,0.0249673782184485,0.00864478558434523,-0.00190149975607645,-0.0230460047360466,0.00539682539682551,-0.00199870871444952
"2388",0.0180363265820911,0.0322489286725753,0.0150709211827997,0.029475692499654,0.0020833462679557,-0.000176549009045179,0.0217168887160057,0.035897577330821,-0.0107357120303128,0.0160213488817786
"2389",0.0170274737925631,0.0221178949190379,0.0131006141879371,0.0253166512146217,-0.00767235012463807,-0.00406510718253994,0.012803325283995,0.0175741186349212,0.00414934567507186,0.014454602712451
"2390",0.013645364275898,0.0221801682772849,-0.0086207122350237,0.00999403054239645,0.00368507886578362,0.00221814597683512,0.0111681571380429,0.00827051413379998,0.00500639717121421,-0.00582893627845582
"2391",0.00210067213327991,0,-0.00173913970580819,0.00960404531580505,0.0138846688944085,0.00264218336064892,-0.000728252228368143,0.000482582469987003,0.0153396298304764,0.0123778149562057
"2392",-0.0071934519708432,-0.028314366932273,0,-0.0213316748755561,0.012520186901066,0.00548243102481361,0.00765208646606497,-0.021702305375958,0.00825478519570799,-0.0283139731648793
"2393",0.00599805932724795,-0.00408503242311342,0,-0.00265102044857735,0.00161577515925915,0.000175766457900517,-0.00361601792151711,-0.0014789891805379,0.00587004706982275,0.0039734554960511
"2394",-0.00062023521052823,-0.00519549018958765,0.000870955972198884,-0.00265803448863222,-0.0000693209669574424,-0.00131870826792879,-0.00883143352670568,-0.00271540505645995,-0.00376250491476637,-0.0283641363814513
"2395",0.0148905445106349,0.0156680887281757,0.00696259079676498,0.0216169632081473,0.00736533132744754,0.00193695222975276,0.0147687366937586,0.01683156070865,0.0060120161086783,0.0101833702572474
"2396",0.00352696864546043,0.0135319938302347,0.0242005807484957,0.00956519991812832,-0.0087743864539982,-0.00527281704007643,0.00721670021425713,0.0131452083361203,-0.00942392707864148,-0.00403234117737061
"2397",0.00726313420749269,0.0149530117023309,0.00590712541316196,0.0140684205504991,-0.0164396937566416,-0.00591839080852996,0.00119418169611518,0.00937006929659256,-0.0165518687900309,0.0188934773809963
"2398",-0.000139440596135576,0.000263147944253861,-0.00167801936960821,-0.00169892974135266,0.0117854315847172,0.00257677010579993,0.00417465064501532,-0.0021420833352106,0.00920176941876893,-0.0125828817108378
"2399",0.00558342299298054,0.0105206107935278,0.00168083985143608,0.0144641501846028,-0.0145425641312551,-0.00416584235600959,-0.00736426033295301,0.00620223766322048,-0.00771512582601408,0.00402422820351811
"2400",-0.00134169942622075,-0.00598644247366897,-0.00335561015515928,-0.00223663940723229,-0.00859644747027832,-0.00382712364613247,0.000837521440999911,-0.0111425923787148,-0.00384831534048036,-0.00267204288248979
"2401",0.00268715552296706,0.00235669904313673,0.00252529996311268,0.00896590244482254,-0.000939358875267304,-0.000267900315262914,0.00251089435268126,0.00311691976122308,0.00157682912572787,-0.00468862042717499
"2402",-0.00101647489932166,-0.00940445642918897,-0.00671723809286873,-0.0102747897571208,0.00564081198281818,0.00268130129216426,0.00453162503677951,-0.00286809910742336,0.00133814545546174,-0.00605644537272443
"2403",0.00416296977667807,0.00870242230759932,0.00845329087557922,0.00505074947777295,-0.00546524408479199,-0.00205058006609582,-0.000237341658139045,0.0105461949476811,-0.0143070514449103,-0.00677045791683872
"2404",-0.00377709673601201,-0.00235279720696102,-0.00754408038454579,-0.00307110926237653,0.00202460232747104,0.00223323960218424,0.00142512260758565,-0.00189741970055002,0.0152325067009531,-0.00545330161916657
"2405",0.00448498969714528,0.00183435398368825,0.00168910740442163,0.00728078337810678,0.00173210679284486,-0.00080215547406437,0.00830069038789816,-0.000712850131790344,-0.00746272566859252,-0.0020562452815841
"2406",-0.00271588387805932,-0.000261516253098781,-0.00337267696147991,-0.0100082429439671,-0.00072041937330114,-0.000803080014592505,-0.000940736380777074,0.00356722784420715,-0.0069647567386586,-0.0109890024443174
"2407",0.000461646135092586,0.00340142254970166,0.000845971418545588,0.00786285508421369,0.00158626960066455,0.000624955205766442,-0.00459109175992511,0.00545016871064874,0.00422410931518202,-0.00416660978580086
"2408",-0.00106114881220254,0.00651864743448805,0.00169071726964698,0.00334346605366731,0.0124532277821336,0.00428207813281101,-0.00709560867113879,-0.00023577968394406,0.0161111031746033,-0.00976298245846985
"2409",0.0011544633486622,-0.000517902787280811,0,0.000277632498434155,-0.00184852216032383,0.000533179856878174,0.00738453223226054,0.00495072553354281,-0.00288990863774041,-0.00281693550467965
"2410",0.00161467358874812,0.00959047030386095,0.0177216031425163,0.00527502206965069,0.00833368781907962,0.00381726915361735,0.00969504424350598,0.00680237718361321,0.010339902543008,0.00847467913859545
"2411",-0.000829054849506683,-0.0107832379688467,0.00331665570894923,-0.0019329974570037,-0.0108417129447045,-0.00347177518895758,0.00351281192252695,-0.00582467401828357,0.00186079242861803,-0.0175070513551416
"2412",-0.00640718378642158,-0.00259526661875809,-0.0123966611581061,-0.00719436812610819,-0.0103027167110172,-0.00239946777416511,-0.0151689176655798,-0.000937202363453293,0.00812570029309945,-0.0014254239409307
"2413",0.00292260420287782,-0.00416356410640073,-0.00502085744441427,0.00334461269404662,0.000578073666931855,0.000534443958742248,-0.00426543752102271,-0.00821023437279433,-0.00475942259125139,0.0164167665089441
"2414",0.0010639519647313,0.00418097185072819,0.0142977258558081,0.00555544602154368,0.00751393751692309,0.00240403144881918,-0.00238004534517533,0.0070952739102188,0.00169688399677059,0.0042135701416901
"2415",0.00817896651514638,0.0033828356220873,0.00331665570894923,0.0116020098593139,-0.0103978207245804,-0.00621788153521508,0.00131181310181239,0.00234860227799483,-0.0178639569517192,0.00419567454347969
"2416",-0.000595785089910428,0.00103711259288142,0.00413222038603522,0.00710021990507825,0.00188388481786728,-0.000536288983060684,0.000953381198474101,0.0023429769322274,-0.000862414719033699,0.00557102644813079
"2417",0.000596140261389655,0.0095853871074818,0.00905355799405094,0.00677869062900394,0.00983644237750081,0.00357722026645813,0.00368877245683241,-0.00233750022312551,0.00408032793345359,-0.00277004539170966
"2418",-0.00247501098308101,0.00384932111169611,0.00326255054249192,0.000269287542103092,0.00386759684973037,0.0026733592703192,-0.00130425780125265,0.00421740129612913,0.00468895752335863,-0.0118056088131202
"2419",0.00464078515582234,0.00792431510737801,0.00731714578915388,0.0129241027233453,-0.00891777048925324,-0.004799022191178,-0.00949757398247675,0.000233261940580931,-0.0069228376932613,0.0154603742383221
"2420",-0.00086912491652924,-0.000760672094613501,-0.00484270612637083,-0.00372133123006146,0.008422114175614,0.00357196319984854,0.00275671977375236,-0.00186587347886424,-0.00211479599145925,0.00761242387006322
"2421",0.00288405321860519,0.00203023089434162,0.0056773392008076,0.0104053164954354,-0.00942310640013466,-0.00293643690108047,-0.000717085371288118,0.00397276300770999,0.00345364201799625,0.0164835036664763
"2422",-0.00515768098523539,0.000506586188822489,-0.00887093916818116,-0.00448890012924796,-0.00266627197608438,-0.00169573290018132,-0.0117226002268247,-0.00256054658052618,0.00492807430938913,0.00810813667656118
"2423",0.00188089728709095,-0.00151876183559152,0.00813663027990819,-0.00636618003763645,0.00599718832910145,0.00160906733814281,0.00290501256219167,-0.000233468686682725,0.000233509767000095,0.0040214617765566
"2424",0.00224388994276636,0.00760664003249811,-0.00484270612637083,0.00934338949735292,0.00158073532964131,0.00178513191310681,-0.00289659790887875,0.00373496968586018,0.00474708949416347,0.0126835420999869
"2425",-0.00146192619821328,-0.00830417980004916,-0.002433070604973,-0.00555406342365761,-0.00523538217253205,-0.00338557062272815,-0.00726222061225068,-0.00697674362126943,-0.00882968004934037,-0.00329593395865624
"2426",-0.0000459693694260244,0,0.0056911206782877,-0.0132978020999762,0.00843492963455916,0.00223492065508757,0.00512074808162999,-0.00210768231034719,-0.00148473859900955,-0.00925926871340432
"2427",0.00201345217566851,0.00456737310909472,0.000808444391098284,-0.00404296541604376,0.00107243661403622,-0.0000895685050313899,0.00218341745833261,0.00657112445725039,-0.000156495540432733,0.00400528569093561
"2428",-0.00511470404082814,-0.00303118472987984,-0.00080779133672304,0.00270602287775157,-0.00235675091917176,-0.000356305860495509,-0.00484126850369293,-0.00373049349893628,-0.0111146366450433,-0.0119681274213354
"2429",-0.000688617219754772,-0.00430693118418468,-0.00485036203606171,0.00080990457428598,-0.0037936780728649,-0.00160648532454177,0.00364856207028574,0.000468340348255714,-0.000870611077112948,0.00403776877017403
"2430",-0.00188329410016763,-0.00534348793597073,-0.00731128802201131,-0.00863012837058852,-0.00582041720670101,-0.00384336887773573,-0.00933126273365403,-0.0112283417270046,-0.00142596843636289,-0.00335122964418233
"2431",0.00492421799637932,0.00460467637374884,0.00327342829729926,0.00761699392777615,0.013371455763092,0.00412789152796877,0.00941915534692539,0.000709893042637466,0.00198333989726285,-0.00403491472006745
"2432",-0.00164862383894904,-0.00152799969006889,0,-0.00269968654071073,-0.00385185504433461,-0.0000898737281379569,-0.00169645564093313,-0.00520102695448466,-0.0100554550263946,-0.00945308182100768
"2433",-0.00284398027309085,-0.00178511778440982,0.00163133009997352,-0.0110991581282369,0.0014318412629164,-0.00116195830239252,0.00194212339939548,-0.00166378228105213,-0.00199952013116467,-0.0190865205881448
"2434",0.0000459087873880826,0.00562079638478497,0.00732895274844259,0.00766507240522341,0.00110326456453969,0.00156836012286088,-0.0016960587061261,0.00928370757932218,0.00408720952145547,-0.0111189659261556
"2435",0.00450802091990732,0.0149899668007656,0.00727556479055913,0.0162998364360423,-0.0081564500977388,-0.00259421619365607,0.00800956070663017,0.00117954799120024,0.0102162901251792,0.0112439874393682
"2436",0.00302242352942961,0.00550657962896084,0.00561795437259804,0.0213847371590923,0.00728568391947126,0.0046633733758481,0.00710326737455591,0.014840723231877,0.0169076953464486,0.00694917489634173
"2437",-0.0000912801815784459,-0.000248886434999318,0.00478859831548006,-0.00314077715045746,-0.000716136746040208,0.000535754762156504,0.00573855535447554,-0.00580301011378648,-0.00341856092044179,0.00897172432975935
"2438",-0.00228305402263262,0,-0.00476577692412916,-0.0026250349356991,-0.0125417815238433,-0.0049071253102555,-0.0114111111542728,-0.00256822668346912,-0.00530137973645028,0.0177838964431223
"2439",-0.0239348010054349,-0.0209162468706494,-0.0159616510423997,-0.0336935002843118,-0.016473901441887,-0.00475210640249057,-0.0397981454476526,-0.0255150099050973,-0.00658355691146817,-0.0154570542315235
"2440",0.0143471132451405,0.00890121774374664,0.00811038799879671,0.006810444348611,0.00051644554186514,0.000901058212525729,0.0121462549578233,0.0048039547903731,-0.001262358974359,0
"2441",-0.0143754572986164,-0.01991403318586,-0.017699145290123,-0.0251625982233958,-0.0113574341705852,-0.00369026216933455,-0.0243721342660431,-0.0207983925238253,-0.00663556384028952,-0.0129693172763443
"2442",-0.00037505231198609,-0.000514605750904784,-0.00655201995235644,0.00305330234156775,0.0014918028526596,0.00225890974876286,0.00304338894287803,-0.00170886212097188,0.00341948310139162,-0.00760708883651384
"2443",0.00999282579623584,0.00797733448666538,0.00494632982544174,0.0171553481603854,-0.00432086206723703,0.000269963291544828,0.0045512396222398,0.00611396854151036,-0.00641937708036144,0.00487798195622902
"2444",-0.00386548434299006,-0.0178706962515262,-0.00820338030618317,-0.00680073002925285,0.00808050917055581,0.00108112139001326,-0.00100691535659447,-0.0110591936192251,-0.00247272068741999,0.00138694364428016
"2445",0.000187472758285789,0.00779808795875048,0.00330853742812165,0.00794288946584465,-0.00326565008630142,-0.00171031314522652,0.00944819560487131,0.00793480518959688,0.002079018104574,-0.00069244007257252
"2446",0.0000469902720583448,0.00206356932554597,0.0140148154486137,0.000543464637077218,0.00349961861751047,0.00153330030151078,-0.00162215223183371,0.00442791852846347,0.000957564634535668,0.00346495601403118
"2447",0.0112453424593375,0.0128701998973748,0.0292683864150753,0.027974214148669,0.00808732136184354,0.00162041657489564,0.0114998759152618,0.00857201449566247,0.0145886078668909,0.0124309117376125
"2448",0.00630155383670905,0.0116899151885528,0.0126380859034478,0.0071331533311445,0.00794860755804394,0.00296630119308672,0.0194021663868242,0.0114133438810065,0.00235721699592717,0.00545709200812983
"2449",-0.00547926263833631,-0.00753583021772342,-0.0140404290412256,-0.0128540249768534,-0.000949401887926471,0.000447930259534823,0.00254557299247926,-0.00408155035660684,0.000627122364192267,-0.0115332945108013
"2450",-0.0081022717182897,-0.0111364887049294,-0.00870267402093405,-0.0146159811864131,0.00635831220198169,0.00286645272465957,0.00117065580943754,0,-0.000783384241545115,0.00686346568920571
"2451",0.00620797195338074,0.000767910799325477,0.0111732887749116,0.0142932971484682,0.00733542549299027,0.0016974645875274,-0.0077952324155045,0.00771450597455203,-0.0072912581585749,-0.00954336553088786
"2452",0.00496351648570159,0.0112532652988846,-0.00157868904337599,0.00904027378173788,-0.00216289969523442,-0.000446127510668193,0.00552402237722838,0.00334928751024943,-0.00315907432098228,0.0233998982825621
"2453",-0.00904730752223459,-0.0144161350798495,-0.00711444086981461,-0.0173914758218325,0.00252898016097869,0.000624581276253977,-0.0107437296158176,-0.0164520161740668,-0.00118840911750584,0.00605251050862865
"2454",0.00754617199977692,0.0105210420120483,-0.00159236524414053,0.00429082359127775,-0.00893665141013189,-0.00249633166985808,-0.00481266792372814,0.0111513704686619,-0.00341081145395405,0.00334226902923129
"2455",-0.0024040971713446,-0.00152353231344371,-0.00318963829624375,0.00694262143591207,-0.00330042174466727,-0.00232686131912918,-0.0181052592904031,-0.00455522565842004,-0.00254695162804008,0.0086608425336514
"2456",-0.00509781224876604,0.0015258570058978,-0.00560014757857807,-0.0111377870822994,-0.0116950723345972,-0.00457534979865515,-0.0143975250373121,-0.0139690513441701,-0.0347111315033514,-0.0026419718257199
"2457",0.00442526455103631,0.00253936297517066,0.00643598990464511,0.014481145392407,-0.00465968853943277,-0.0022531378739391,-0.0193490786693963,-0.0134345125903319,-0.0015706538681437,0.00596018324407677
"2458",0.0006955903752075,-0.00607894901070483,-0.00479610312564205,0.000793088921402507,-0.00557284796892465,-0.00207724978969948,0.0016988183688762,-0.0118839988847488,-0.00927301713258011,0.0019750244006882
"2459",-0.00342927127677506,-0.00764529661904412,0,-0.0044902888809667,0.000672870225327582,0.00144836886922439,-0.00143528514852453,-0.00876974562582644,0.000668510758197849,-0.00262808499404299
"2460",0.00520831972584213,0.00231153872927292,0.00321269587401241,0.0108781780387428,-0.00589910332593424,-0.00262162023066514,0.00587868893468246,0,0.00350764996672215,0.011198928205062
"2461",-0.0126295202964029,-0.0148606632439534,-0.00880686822744725,-0.0230971706554625,-0.00225344706367936,-0.000271787011396296,-0.00999997429787769,-0.0171890930083848,-0.00507657273380246,-0.00586324608441957
"2462",0.00131191990137047,-0.00286059881273215,-0.00161575642470813,-0.00188054384663561,0.000978616828528622,0,0.0135117642659528,-0.00154312200135476,0.00158925131938314,-0.00720842462624149
"2463",-0.00327546956833635,-0.00443422008273164,-0.00161795799148023,-0.00888300999883018,0.00376043427486561,0.00208519062841628,0.00556558659500417,0.0108190816621758,0.00242192253920037,0.00660070625287879
"2464",0.000516432784268384,0.00104797391367106,0,0.00162968793080531,-0.014011462377879,-0.00307553556787232,-0.00334657859309062,-0.002803129815937,-0.00558192123287449,0.000655728765314612
"2465",-0.00347230117460451,-0.00366411289368296,0.000810497009395172,-0.00108472079743305,0.00638316039730502,0.00217752769113466,0.00129146646081657,-0.0053668002414492,0.00268095674697588,0.00131066557908799
"2466",0.00626241723773613,0.0123459293332666,0.0056678176402698,0.0176438717791692,0.00324712312444442,0.0019916289360038,0.00683588563196658,0.0125899805581686,0.00618313836898388,0.00196339129656375
"2467",0.00266710304339268,0.00155659263705776,0.00322062962588276,0.00613493307321678,0.000828151481389261,0.000452042727496327,0.00422771243051079,0.00558223987559692,0.00572997019980015,0.00653165629159558
"2468",-0.00186665959663435,0.000259242056333875,0.00882830958027836,-0.00291618100904167,0.00105289490117433,-0.000903306195120246,-0.00382705507185055,0.002523806656761,-0.00305509864540421,-0.00908501892228064
"2469",0.000467440014894738,-0.00259000514891738,0,-0.000265850758030761,0.00150273317164862,0.00108495333330549,-0.00128066988056097,-0.00226576314927696,0.000745436487418205,0.00392921932243606
"2470",0.00425280749489598,-0.00129842361578125,0.00159109852429951,0.00425532950180152,-0.00435126001987418,-0.00135490964155571,0.00269277972559379,0.00227090849004918,-0.00223457746859923,0.000652373967855002
"2471",-0.00335082687764765,-0.00260001921856068,0.000794317510661502,0.00105944135272473,0.00263696431529126,-0.000180430192231573,-0.00191795478618395,0.00125792861587293,0.0075481338345742,-0.00456323801298775
"2472",-0.00200748677183304,-0.00547442859050262,-0.00158731012317737,-0.0105819183279048,-0.00676313035510778,-0.00217089726000763,-0.0116593673997686,-0.0103067784156486,-0.00559809001730394,-0.00654883367309145
"2473",-0.00266680496044003,0.00183483470297952,0.00158983368227528,-0.00855628651954921,-0.0108938343944334,-0.0034439774074424,-0.0229453855127262,-0.0111755960905677,0.00182135109014525,0.0059327489710721
"2474",-0.00295536553243037,-0.00130830492698863,0.00158739548193543,-0.00404550271356763,-0.00221803991592551,0.000181558987158104,0.00199021615640183,-0.00616515704754228,0.00471035443830492,-0.00655305811402018
"2475",0.0000470295246925989,-0.0010477093702882,0.000792194808079349,0.00568653033251421,0.00613278401394557,0.000818561663735951,0.0148304546421276,0.00749557953344882,0.00296101327585108,-0.0131925678921104
"2476",-0.00724532911265929,-0.00445861190156049,-0.00395873279930992,-0.00807757903978079,0.0000760437165796546,0.0000361695065422829,-0.0220509044544919,-0.00384828944830296,0.00647860412533041,0.00467914912177814
"2477",-0.00601868876301681,-0.00711284608009632,-0.00635914236655744,-0.0119433598687481,0.00435111643678665,0.00300293214651659,-0.0128086554652486,0.000772704509771183,0.00741461727170334,-0.011976089318696
"2478",-0.00457715461776731,-0.0021224919670908,0.00239972215441675,-0.00274736504450324,-0.00767614542209716,-0.000635192674426244,-0.00581177725844462,0.00257318242977034,0.0053381106869792,-0.00336702670285538
"2479",-0.00110175174693905,-0.00904009840295084,-0.0119711095283497,-0.0101928241162856,0.00896062485525451,0.00308601729142199,0.00530181720016998,-0.00769986731696304,0.000724022508671984,-0.00675673420271494
"2480",0.022057107769609,0.0160984835086506,0.00706770181008198,0.0361813514181808,-0.00850195274173293,-0.00416222786413123,0.0163624620145226,0.00931168565843099,-0.0180078544738954,0.00408164694177549
"2481",0.00450392930599919,0.00316888712841235,-0.00120310778185984,0.00644643035557668,-0.00405713940834196,-0.00354415846750555,0.00612038860497921,0.00256283036433347,-0.0041752189246792,-0.00135499503103398
"2482",0.0106021020839162,0.00500138051911958,-0.00843183417888682,-0.0325594767103103,-0.0424324427325461,-0.0152289421329553,-0.0185133874518252,-0.00434571408479856,-0.000657686621651554,0.00474898719275374
"2483",0.00249560297461371,-0.00366684494178637,0.000809830363741382,-0.0284137223314028,-0.0147703723939708,-0.00601882350299243,-0.0181894751378493,-0.0269576171011647,-0.0148897501627139,-0.00810266141648341
"2484",-0.00230506578172962,-0.00972649535239889,0.00141601829381011,-0.0190232753845252,-0.00562226902028651,-0.00204983254635682,0.00535213024506942,-0.00765178633065577,-0.0221294530271399,-0.0190606052729353
"2485",0.000785654550988113,-0.00822957607363106,0.00121218755398655,-0.00723580451703454,-0.0059817984403977,-0.00578758264526025,0.0169256523776566,-0.0124964425828747,-0.0084542870786386,-0.00208185917709702
"2486",0.00780261024699613,0.00588880766172339,0.00161412686856188,0.0201166267131585,0.00494600399326717,0,-0.00362392608661621,0.00700049925425428,0.00869866498407834,0.0222531114282418
"2487",-0.00187832534556076,-0.0119744659370578,-0.00483466365070295,-0.00828806297243301,0.00902339004657082,0.000938950082886469,-0.00215541256784646,-0.0131015898839957,-0.00298843913110214,-0.0122448708106266
"2488",0.0051408217490081,0.00457848215520573,0.014979558909979,0.00144098122919312,-0.0147146076311764,-0.00440907843651483,-0.00823572564456232,0.0149010734736781,-0.00513829763993223,0.00206601655464245
"2489",-0.00223762773828917,-0.0109920883325502,-0.014957885779854,-0.00460461276386825,-0.00288751029650591,-0.00442830972907149,0.00299508103793844,-0.00854238461867152,-0.00878020158010162,0.0082475228783081
"2490",0.00755141330991815,0.00975890525614043,0.00809873915886383,0.00982969536126821,0.00248228266767203,0.000851780320721751,0.00013571495060094,0.00215403997030261,0.00373425959645224,0.0279482321863713
"2491",0.00195348363381842,0.00107385665801196,0.00240999494684768,0.0151732001354126,-0.000330284545470239,0.000945527577743244,0.0170988156299665,0.00537326440100738,-0.000346089282815432,-0.00132631000327676
"2492",0.000543798605181056,-0.00724055381687372,0,-0.0107162167521589,-0.00388061920608673,-0.00358984308433186,-0.00547038209104789,-0.00213771495799142,-0.0198199842494375,0.00398407763104802
"2493",0.00371538969316032,0.00810367471468809,-0.00841502616040224,0.00484584946857081,0.00149212629801276,-0.000853468160635029,0.00509783804068986,0.0013392416552358,-0.00565120529801322,-0.00727510080633487
"2494",-0.00469467164778181,-0.0112540905839031,0.00868856978575083,0.00397168807076587,0.00736643722296049,0.00455501882948806,0.00347041885594401,0.00748819309840676,0.0105674628312986,0.00333106690960094
"2495",0.00195040699479088,0.00840106254580752,0.00100159987962445,0.00141266844788945,0.0041901799612527,0.00103909233994504,0.00824659697215391,0.00398218601130895,-0.00465734609866397,-0.0199203198141998
"2496",-0.00239925352411074,-0.000805934237707917,-0.00160103377372844,0.00169311552600293,-0.016200232557991,-0.00670012439734624,-0.0125325740565567,0.000264400983798874,-0.0134192375762137,0.0304878065787826
"2497",-0.00367549653131927,-0.00134499115047682,-0.00841839965619573,-0.0118307826365619,-0.0105587030617302,-0.00381498752477982,-0.0157650881446719,-0.0129526682818182,-0.00187918568232659,0.0184088928598929
"2498",0.00050077631467671,0.00296262726311491,0.00303200197963571,0.00114006496237007,0.00732752620798172,0.00448852155222301,0.0105876121108235,0.00723059504786572,0.00537921816945297,0.00710139187360448
"2499",0.00600881604324877,0.015843223824356,-0.00120908267273467,0.00825744719744992,-0.00108708289872361,-0.000380310344220147,0.00792505327527859,0.00452012163201365,-0.00535043700151983,0.00512820106818124
"2500",0.00316750245746134,0.00978036855849362,0.0044389736714745,0.00536589237525775,-0.000753591429982325,0.000380455035205562,0.00639646977128461,0.00608814191558205,-0.00098620225043744,-0.00446429040277008
"2501",0.0130806432318746,0.0141363172401199,0.014865386345069,0.0168537539607891,0.00854452238233039,0.00332770783054426,0.0194649611818281,0.0142065551139581,0.0035897155164677,-0.0076874068323729
"2502",0.00244884963401382,-0.0043883200438497,0.0114806487108541,0.00442002205200565,-0.0117939366135121,-0.00379033668150586,0.00506555441487766,-0.000778115506416821,-0.00232497536752252,0.00193683988393856
"2503",0.00604027416268527,0.00518517874253877,0.00293537092604823,-0.00522581497612262,-0.0124391046140463,-0.00513657443266158,-0.000775368733517912,0.000778721441645702,-0.0104866720444563,0.0051545684159735
"2504",-0.0011477606865844,-0.00154735866714761,-0.00975605139229219,-0.00663513708693986,0.00187230818243456,0.000190954900984197,0.0062081822853417,-0.00544724489646586,0.00380432964122579,0.00641030081676885
"2505",0.00667399111943068,0.0116246823752348,0.0118225654525168,0.0111327848627745,0.00356774697477324,0.000573671823428157,0,0.00808529674364378,-0.00333877458942422,0.00254773579355727
"2506",-0.00825411761214478,-0.0145556001963942,-0.0153844465365138,-0.029727629178851,-0.0111732527174829,-0.00831155282418561,-0.0185089811231522,-0.0165586120604729,-0.0146672253870682,-0.00952992615734338
"2507",0.004117045058327,-0.000258960334295177,0,0.00170230389612325,0.00505072521768968,-0.00279402849237387,-0.00746479614197915,-0.0144700088905011,-0.013691132708056,-0.00128285619031576
"2508",-0.00195573402114868,0.00311033555726015,-0.00870267402093405,-0.00453117996991714,-0.0023000288026741,0.00125602027557603,0.0133264561357922,0.000739237183633668,0.00661456145386863,0.00449589628991709
"2509",0.00217736149478953,-0.00361748775667137,0.00857950760517667,-0.00682802108075709,0.0107567918354006,0.00463152625074792,0.0110676715913232,0,0.00499762133278225,-0.00575452855061109
"2510",0.00385765964753193,0.00363062148544402,0.000988968118299294,0.00343722917017431,-0.0049833240892414,-0.00211315122686062,0.00180304656920871,0.00653393536837599,-0.00736711510699384,0.00450167871434171
"2511",-0.00278256642237362,0.001550389170063,-0.00533808903295097,-0.00415746981280918,0.00441375791514043,0.0016361353608958,-0.0123057250459171,0.00028229666581292,0.000556610069982311,-0.00576196249489347
"2512",-0.00172776239427541,-0.00179356942749442,-0.00160794190167957,-0.0118876036191161,-0.00178754347629373,-0.000433006448589346,-0.00184750129328848,-0.00395048942982157,-0.00241077426816461,-0.00128774623731354
"2513",0.00146452171483702,0.00286448017040319,0.00181196303129671,0.00586833954508759,0.00203692916548182,0.000962860498859186,0.00264431927333186,0.0048160633792218,0.00316018229055426,0.00193420953618118
"2514",0.00248091351434399,0.00129850670138998,-0.0062298986250604,0.00437593489790356,-0.0032185910890673,-0.00144317042120534,0.00118667292940344,0.00535642285192872,0.00583709811915112,0.015444003425422
"2515",-0.00826451404666084,-0.00622429879175468,-0.00141560553045217,0.00755145141948543,0.00730833007014642,0.00366079898973792,-0.00592702356742636,-0.00701043345287511,0.00276347646948194,0.000633704922959666
"2516",-0.000222817638010131,0.00704609931478983,-0.0101254915758263,0.0164312081567819,0.00354326875199518,0.00307149797065231,0.00993755334947877,0.0104489878211058,0.0131361380384334,0.00126673755373652
"2517",-0.00365493331290168,0.00570101333072959,-0.00040920004544831,-0.00709014903705085,0.00151354344235632,0.00296623062654855,0.00944642608061996,0.008384698326249,-0.00616556345846808,0.0018974420434541
"2518",0.0076500199399907,0.0023189402779773,0.00818656786143079,0.0119965808625599,0.00428108263174876,-0.000477215913189388,0.00402915922530744,0.000831430623377871,0.00784599938102359,-0.0119949157764663
"2519",0.00594937811162555,0.00874021445870876,0.0200975971870214,0.00762071629197059,0.00384468040167785,0.00114528398253855,0.0137217837685066,0.0105234458930408,0.00353037020430547,0.00766769250680732
"2520",-0.000794605475076704,0.00866476877699074,0.00577102059246903,0.0109242524766051,0.01565361108003,0.00648299333971725,0.00344772785644087,0.0150725587353084,0.0155150729251752,0.00507298460463712
"2521",0.00357765615817485,-0.00429512555241018,-0.00158297607706281,-0.00415622951935346,-0.00918175046514513,-0.00454656344439275,-0.00216329967711504,-0.000270026178959326,-0.00737255272033122,-0.00126187729913718
"2522",-0.00330081547590799,-0.00380619121185966,0.000990968168421258,-0.000834727299524163,0.00802567454083203,0.00380618945480138,-0.00663200390683849,-0.00189052973516601,0.00823264429530202,-0.0151611396094232
"2523",0,0,-0.00376163534801488,0.00584791186926892,-0.00065630305860942,-0.000473716049096629,-0.00937212004888721,-0.000540925563579986,0.00426026456483997,-0.00448993064839287
"2524",0.00282614251772317,0.00534902144399108,0.00655803670755439,0.0119048017702121,0.00336728738654379,0.00113784292424679,-0.00427679463640751,-0.00243632116655024,0.00309322133286405,0.0109535241994081
"2525",-0.0025101357307209,0.00177347352826529,-0.00157943324692711,0.00437757946616157,-0.00221035767664657,0.000568310515377757,0.00455526692553043,-0.00407078191786148,0.0036123700440529,0.0146590152638848
"2526",0.00229580596142931,0.00379359273297419,0.00632779027916697,-0.000817099975730651,-0.00475836375441874,-0.00217764606715454,-0.00103628467779404,-0.00108994580529775,0.00263361416438879,-0.00188439640516536
"2527",-0.00352364751819689,-0.000755710876173765,-0.0112005992794416,-0.000545317419389124,0.0104693629842929,0.00502864730416208,0.00674458470077455,0.000272891482451687,0.0143595045474083,-0.000629382790976241
"2528",0.00220993316095375,-0.00378231049946898,-0.000198660521451455,-0.00545567394221624,-0.0128082491525866,-0.00708054188488649,0.00167457062807186,0.00054533586911143,-0.00845917148828956,-0.008816065726727
"2529",-0.00370433838274509,-0.00253094468957782,-0.00278283538025526,-0.00301683580335932,-0.00685873170588636,-0.00380329488876474,-0.0104179038813805,-0.00981178831254226,-0.000870601526840709,-0.00317664205244783
"2530",0.00367397665006863,0.00532846425971267,0.00637847456502572,0.00192551847984523,-0.00199725152397001,0.000477443756947915,0.00636860643327708,0.00385364457859128,0.00243971427480294,0.0114722499988849
"2531",-0.00260221518816084,0.00328147003427004,0.000594059034850769,0.0148270986149459,0.010005193702066,0.0052470048183324,0.00761990465998652,0.00795168198175999,0.00643196854153927,0
"2532",0.00641178067668213,0.00201245752076984,0.00257322550028594,0.00622296445503312,-0.00685165026373824,-0.00379638143350192,0.00230717990612561,0.00108816657928856,-0.00449092318429123,0.00252050941723025
"2533",0.0086553660449753,0.012051025203675,0.0104639551579322,0.011024446843827,-0.0125507753722329,-0.00495347954499081,-0.00537106190869696,0.000543376324157796,-0.00824149409841668,-0.00628526933019513
"2534",-0.00104519626301136,-0.00620184346189867,0.00136769261684866,-0.00425530435014476,0.00336680289052049,0.00134024592057669,-0.00102862802131876,-0.00461698237896435,-0.009272200839748,0.00442745156679414
"2535",-0.00157000837021526,-0.000499200345479123,-0.00819498901980076,0.000801372024345381,0.00360757481590857,0.00124304372913286,-0.0093951556154952,-0.00136446474851504,0.00203069041090065,-0.00818635137568224
"2536",-0.00620160833509387,-0.00874130089466252,-0.00275436638738935,-0.0053376206461051,-0.00300933081294741,-0.000286711843741183,-0.00688539936784349,-0.00109272464218724,0.00422947403699836,-0.00571427301828686
"2537",-0.0000879178944857006,0.00377914355254982,-0.00236730131320595,0.00187830925443944,0.00695892854962854,0.00343877556314398,0.00784902932650877,0.00957337020476579,0.0138633147857918,0.00574711359443247
"2538",0.000395603705494851,0.00326323785575044,0.00533904085671888,0.000535474398245084,-0.00618316767777793,-0.00191631536044223,-0.0118120533729819,0.00189641263616291,-0.00302904362538192,0.0107936340731034
"2539",0.000658991929602504,-0.00100078802689452,-0.000393173551912374,0.00428266923648613,-0.00041983021833536,0.000382312533736329,0.0111652829205431,-0.00243358740945254,0.00555554701967576,0
"2540",0.00689290491545202,0.00400696721760663,0.0045257009393207,0.00612996773465802,-0.000419878180312305,0.000763461263792564,0.00675487540345676,0.00542136251197944,0.00250346175771621,-0.000628132135055082
"2541",-0.00178788770677318,-0.00947865363482236,-0.00156716166453474,-0.00238408507747534,0.00605042936891698,0.00477069002608377,-0.00335478396723743,-0.00188747146632151,0.0135193321325926,-0.00628526933019513
"2542",0.0000437693255843641,-0.00125895857575919,-0.00058863153336719,-0.00504504178140885,0.00735051178403312,0.00180419695216605,-0.00142407231605124,0.00216111441405342,-0.00203906547253352,-0.00442764686394759
"2543",0.00131052143714139,0.00252125956285476,0.0029446615502926,0.00613806017243945,0.0135985054184755,0.00407564360989454,0.00726049800410089,0.00539084043448312,0.00621490725536278,0.00381195738522355
"2544",0.00593262552183926,0.00402409973213858,-0.00137008113695358,0.00450941481575429,-0.0115344429511459,-0.00594725271360841,0.00308912043556142,0.00428961973977526,-0.00761486576504167,0.0050632218761828
"2545",0.00394607381732959,0,0.00705605160461453,0.00924214571988147,-0.00057952388392668,-0.000664646032312866,0.00769916435225748,0.00106770274602863,0.00264299597030426,0.0107053384040592
"2546",0.00544272571308757,0.00450903391170177,0.00389258553756267,0.00313978474144916,-0.00314688901054527,-0.00152021882154052,0.00331100056808209,-0.00293294562619995,-0.00680267868712037,-0.0112149924655612
"2547",0.00399530674223292,0.000748289655380763,-0.00717341700677809,0.00104332859024159,-0.00722684268705764,-0.00361688049683706,-0.00558459022139801,0.000267173501275808,0.00111298798511172,0.00126028713508397
"2548",0.00522022203707895,0.00274099271269024,-0.000976371786166608,0.0080769788344035,-0.00460230671959083,-0.00191020862375413,-0.000893667234029061,0.00187153420193842,0.00444707944924305,0.00125863603933829
"2549",-0.000851280387739295,0.00472178463047945,0.00117280784803331,-0.00361832094823111,0.00546389500249633,0.00401921001233818,0.00472672841365229,0.00080065261034723,0.00536402738264852,-0.00628526933019513
"2550",0.00157643399990115,-0.00321564370602745,-0.000585675478290693,-0.00415055177873758,0.00593609590433064,0.00266914289425135,0.00165297457059999,-0.00106656397274618,-0.0033875507556308,-0.00189763734060744
"2551",0.00595512966443223,0.00124083119636476,0.00840018973074375,0.0109404696042383,-0.00174546052206426,-0.000475358741078624,0.0125665159606358,-0.00240269606376431,0.000594833446634802,-0.00126734462309919
"2552",-0.000888062789811572,0,0.0011622122816124,0.0030919400830407,0.00166516342694734,0.00161682698783761,-0.00250719624930118,0.00240848291618678,0.00135884501061567,-0.00507620312805912
"2553",0.00067703227921756,0.00272604817809463,-0.000967492212295529,0.000256704174791844,0.0029922388951098,0.00265900441021505,0.00427288362699807,0.00453793938462188,0.00873545895223615,0.00318873197427805
"2554",0.00126895117278969,-0.00889768035014182,-0.00213058121625487,-0.0118129731147669,0.0111047838309093,0.00464069883244611,0.00500582202700817,-0.00212582350234125,0.00638973421238043,-0.00190709233946518
"2555",0.00156298756398043,0.00174561117439942,-0.00310554462609047,-0.0031185982287929,-0.00590109385353121,-0.00358229181071568,0.00522972055014925,-0.00399457226108579,-0.00484539694683539,-0.00254780134871879
"2556",-0.00269914022839557,-0.00174256932591199,-0.00253107798291896,-0.0096452975091168,0.00371004117242002,-0.000473146372884981,-0.00396382201611811,0,0.000923438526105436,0.00383143097049166
"2557",0.0139975438572957,0.0117207424215227,0.0117119067624534,0.0155304521842332,-0.0167564205076957,-0.00696644206766739,-0.00310905083817625,0.000801988627725292,-0.00142585755030133,0.00445286527660071
"2558",-0.00629748519693896,-0.00369739012712378,-0.00945404838192176,-0.0176258527985861,-0.00359902780816079,-0.00286334076382688,-0.0041167206510071,-0.0125568220567593,-0.0124306738187582,-0.0158327854283856
"2559",0.000629536840404121,0.00841173164048148,0.000584327220758851,0.00765159636161616,0.00260421209493922,0.000957054225466214,-0.00238019739135198,0.00405860181441997,-0.000595339333299139,0.0051480673719293
"2560",-0.00297786666343713,-0.00515206412035518,-0.00233604740497628,0.000523784680868999,-0.00477603807926252,-0.000191143733831889,-0.00464579538127041,-0.00161680643160456,-0.00672284049488825,-0.00128045807361343
"2561",-0.00298682434238995,-0.00567194088397938,-0.00234137209258722,0.00104687835669304,-0.00303083544792138,-0.00143503169419823,-0.004289053928061,-0.00485843814957099,-0.00805347834087144,-0.00448725015697193
"2562",-0.00185665656124279,-0.00421618585198225,-0.00312931538561245,-0.00941179554047056,-0.00540477749665924,-0.00335234269326989,-0.0153300261562124,-0.00867903284016802,-0.00621869931092334,-0.0225369177448197
"2563",0.00126810215322348,0.0079699934264037,0,-0.00791759628233868,-0.00798053513576158,-0.00278705371046051,-0.0127380082122024,0.000547059808659212,-0.0051277334456411,-0.00856391818071489
"2564",0.00350433947241502,0.00889539834031905,0.00725918403167247,0.0111731916451974,0.00350901427445294,0.00212048311319779,-0.00247636047880917,0.000273729196672345,0.00218397831585593,-0.00930240351013967
"2565",0.000504813018472827,0.00391883421582007,0.00506425207699879,0.0139437728658816,-0.00631120536951257,-0.00250086527475579,0.00156770754775293,0.00191355394184733,0.000174311365286783,-0.00134129435353814
"2566",-0.00382657617830506,-0.00731898227796091,-0.00697673963416223,-0.00570834475842963,0.00480606165888475,0.00106077470953769,-0.00091314529624098,-0.00818579395909336,-0.00540347752141324,-0.00402956400638621
"2567",0.00865352853578094,0.0135169513116966,0.0101482919027203,0.0260958314092532,0.012215290748969,0.00876439432489651,0.0184099152057997,0.0159560035026385,0.0186645368384717,0.00876603378785168
"2568",-0.00196709456979205,0.0104267750038753,-0.00193209644407932,0.00610372902908352,-0.00506344690354465,-0.00276870305712185,-0.00166674909665987,0.0119145041402662,0.00412905806451613,-0.00133694889041081
"2569",-0.00175620022522749,0.00191970436584832,0.00329096555088637,-0.00176916710401409,0.00627647595327741,0.00268082134917846,0.00423801968000515,0.00263645956555147,0.0022273193979101,0.00334674345417874
"2570",-0.00109679389440209,-0.00191602616205988,0.00019287278547564,0.0116484442365825,0.00429883532608488,0.0023869359572164,-0.000384172703450703,0.000804899647445456,0.00444485861090449,-0.000667102292611355
"2571",-0.0128395918016989,-0.00359978640022085,-0.0077161922732667,-0.0110139657141992,0.00830881614030021,0.00333342190204533,-0.00319757391976017,-0.00750680845812146,0.00876520281226778,-0.00534051833327187
"2572",0.0023532377144897,0,0.00136094519245344,0.00480892531773169,0.00399524990768407,0.00189933641230278,0.000513045582033245,0.00270141160337389,0.00244643999960825,-0.000671062731966487
"2573",-0.00106715226519072,0.00120415661593665,0.000776531670744207,0.000251917460224016,-0.00140926047466639,-0.00104273292446067,0.00743965044355055,0.00404092371710152,-0.00134649497018424,-0.00201488568513231
"2574",-0.000726430870895411,0.003608553691691,0.00620749496730855,0.00251848525589304,0.00356973591400278,0.000569296063311908,-0.000707007973123619,0.00295139598789529,0.00160110392855994,0.00336476113458128
"2575",-0.00102620129363862,0.00527308682017891,0.00057850017869443,-0.00276337973856555,0.00455020730529787,0.0024648342839384,-0.00681745186473615,-0.000534923712668722,0.00563686685481346,-0.00134129435353814
"2576",0.00727690104597256,0.000238398339118318,0.00847774263786616,0.00277103716652638,-0.00667066320690635,-0.0034044856962675,0.00440349208051427,-0.000802960583149548,-0.00409937257675375,0.00604431144893303
"2577",0.000934836260128469,-0.000953445708567924,-0.00133738077787215,0.00175824812301162,0.00596927550041926,0.00284691922179259,0.00438430297343961,0.00267858903233753,0.00243616429405091,0.00934580402420737
"2578",0.00318413478138035,-0.00381774137533542,-0.00554813966746681,-0.0052659508468812,-0.00807650934267889,-0.0028388372813688,0.00295296064737594,-0.00534315731477186,-0.0072069134801489,0.00396826774429404
"2579",-0.00232760587299319,0.00239515272425872,-0.00923422654606609,-0.00705819911678707,0.00290803261977324,0.00199284447293113,0.00473609625271831,0.00456622546126551,0.00211023886122863,0.00197625751826047
"2580",-0.00173917877901408,-0.0038231353743805,0.00504845636227258,0.00558524777095371,0.0100865766200597,0.00492274516413627,0.00089185025165972,-0.00106950140172324,0.0053065784593449,-0.00394485458956617
"2581",0.00063735507288798,0.00143920798608055,-0.0034775148006656,0.000505117210659378,-0.00542443324481245,-0.00141571600613222,-0.000891055563531085,0.00214132526797139,0.0022622958066576,0.00990112731437764
"2582",-0.00297262978019353,-0.00670643829651896,-0.00697952694493709,-0.00302832078670645,0.00305760711491976,0.00189029746588831,0.000255053040316255,-0.00160268339233294,0,0.00196069013709699
"2583",0.00281110570621146,0.00337591284240202,-0.00507611705605637,-0.00177159900772794,-0.00148310688935271,-0.000660660924586831,0.00687800911908987,0.00909580465911608,-0.00367833965026731,0.00260929445926572
"2584",-0.00101931909309472,-0.00144226919732182,0.00215859315553013,-0.00177488128547376,-0.00404282944400791,-0.00302053479657982,0.00113856379929445,0,0.00234937909045141,0.00260250376062299
"2585",0.000595079424258627,-0.000962517429967114,-0.00234985324372206,-0.00406399383554756,0.00463940707356958,0.00179908839509557,0.00694979277515029,-0.00397664616298099,0,0.00778704458108392
"2586",-0.00118966087316064,0.00602263632448286,0.00510310083632004,-0.00229531255944682,0.00948274735247279,0.00463130368756093,0.00552130799607387,0.00904986894944892,0.0144818601580603,0.00193185131067319
"2587",-0.00438191580561931,-0.00119734292956897,-0.00331955196802203,0.0048569501090896,0.00547325151085998,0.00310451973092452,-0.00224642205175085,0.00580310799561246,0.00684870852630226,0
"2588",-0.00649495879976469,-0.00695268975859509,-0.00842481379265836,-0.00432464072508698,0.00308686236211853,0.0030018305652697,-0.002001310687191,-0.00209798827418783,0.00475332744025558,0.00321332361178372
"2589",0.00885995723191657,0.00627714055426121,0.0106698944656443,0.0104751950260509,-0.00307736296620353,-0.00158962617645386,0.0125330728691908,0.0113007444535693,-0.00293637851445971,-0.00576545622459146
"2590",-0.00298429926787791,-0.00527836184757269,-0.00312809169799599,-0.0126424035453118,0.0130794914201997,0.00571271222714742,0.00235181223653202,0.000519789289042949,0.00474478083679286,-0.00386605894290903
"2591",-0.0018386103200323,-0.00337672769745556,-0.00058840063258947,-0.00614568067926446,-0.00545300639817226,-0.00260747535236494,-0.00160562590163138,-0.00831139764018973,-0.00887475166910923,-0.0174644522676406
"2592",0.00813912618393897,0.0077444277662797,0.0060832814321059,0.0123678164869743,-0.00387050638456032,-0.00224073749001386,0.00061853081404184,0.00392857545314884,0.00188939451517145,-0.00394991328905014
"2593",-0.00318683665799002,0.000240329845827336,0.00370579157614936,0,0,0.000467656158918084,-0.00395539560258396,-0.00495713260625308,0.00286978519899783,-0.00991407848530956
"2594",0.0109980136784069,0.0362544587157749,0.00699572029828421,0.014252842691971,-0.00493759608313937,-0.00205774088326238,-0.00868699976099019,0.00498182818920867,-0.00678599471483921,-0.00333780678179185
"2595",0.00581848345062874,0.00880442941064108,0.00366648037640593,0.00878302047996926,-0.0120393196295513,-0.0051549447246394,0.00287918291087941,0.00417423993670774,-0.0101251479224939,0.00468855149106728
"2596",-0.000628680006188209,-0.00390448023173395,0.00115366110126369,-0.00373130140999189,0.00551689396203181,0.00263808834810497,-0.00661574784306185,-0.003637485096051,0.00490641164241157,-0.00533332912498308
"2597",0.000838791341773337,0.00069169050932083,0.000768343637771896,-0.00124849794299986,-0.000327726584223975,0.000657439643779512,0.00113086727696698,0.00130403586810846,-0.00372390776974207,-0.00536192604130525
"2598",-0.00217936089796211,-0.00115220027610019,-0.00479766520604008,0.00149997774319721,0.00221180208186533,0.00103293339337829,-0.00928833483242919,-0.00572902641674378,0.00315639175310567,-0.0026954503170562
"2599",0.00252017139531957,0.00392159401232295,0.00385649560861911,0.00574132552351148,-0.00831330967673471,-0.0021608214229375,0.00608151985760563,0,-0.00910821418667418,0.00202706893995463
"2600",0.000377140185202407,0.00689339820354529,0.00307341358082014,0.00719802968609806,0.00512058395287651,0.0020717174533158,-0.00251900174179431,0.0112623911087262,-0.000167092841432237,-0.0107889326307644
"2601",-0.00121455702478235,-0.00251028094537831,0.00248945528995903,-0.00665346460635619,0.000657360797936102,-0.00206743431356471,-0.0119932947948598,-0.00466206938085512,-0.0139573670880507,-0.00408999375384422
"2602",0.00117406435069034,0.0148709726529566,0.00248335452448711,-0.0111635991107464,-0.00492666428476696,-0.00225943491657776,-0.00434441190172652,-0.00208198761826828,-0.0100864720269586,-0.0239561487734999
"2603",0.00393706877081312,0.0114967146219407,0.00552593833899517,0.0082790033506015,0.00090765324958153,0.000188828658449269,0.00962556032500883,0.00573678089575491,0.00188373146773069,0.0140251252850372
"2604",-0.000166956830504827,-0.0104747433907374,0.000378954819640454,-0.000248846030084238,-0.00544167867958656,-0.00245298761531976,-0.00572040179833433,0,-0.00222204935950687,-0.00414932118355293
"2605",-0.000917911952627359,-0.000225189780512114,-0.00322027840956629,0.0126929775788105,-0.0000826898487965577,-0.00113506823565912,-0.00536948521353697,-0.00103690205051354,-0.00599569164882219,-0.00486111622344032
"2606",0.00179583925913263,0.002703111795749,-0.0045609463338333,0.00663537049462515,-0.00116076682081556,-0.000378873768641208,0.0053984722303535,0.00103797833237484,-0.0000861869861390474,0.0160502406843015
"2607",-0.00204284420345602,-0.00292048299135195,-0.00267286065808736,0.00219724632828111,0,0.000758024608834118,-0.00536948521353697,0.000518451025256716,0.00396414164112247,0.0041208935885988
"2608",-0.00167084957600372,0.00788637311844553,0.00248842072161959,0.00414133150510576,0.00755310861667535,0.0051110017336502,-0.00269916346014598,0.00181417070636058,0.00283263519313293,0
"2609",0.00552346571321527,0.00581273481189215,0.00286441797546821,0.0101892357640951,-0.00271846408142384,-0.000659022627114703,0.00360878029884537,0.00517319030481045,0.00265340233410249,0.00547195189069516
"2610",-0.000915601188674509,0.0102244438899186,0.000761456600060884,0.000960853483464863,0.00371695788986193,0.00131930739057151,-0.00565047006845376,0.000257664187834683,0.00435379037351713,0.00136059565705837
"2611",-0.017743961839924,-0.0138613605225542,-0.00152197694661549,-0.0170345749064847,0.0145670001245115,0.00799901286208393,0.00529537561248317,-0.00360220305983294,0.0181895364523665,0.00679338516144568
"2612",0.00402845872215818,0.00133877549073391,0.0026676866865627,-0.0165978275524001,0.00113545702869255,-0.00028018345048364,0.00269745589954429,-0.00335632229531135,-0.00818100836312718,-0.00269901859172683
"2613",0.00650413278147211,0.0131461067236336,0.00817168372918475,0.0213453196998639,0.00234954582069702,-0.000280192079503805,0.00589382915115966,0.00595833480096908,0.00496594571106734,0.0196211203497609
"2614",0.00507733786201148,0.0024191149607844,-0.00056547217708347,0.000971977263914514,-0.00274810613309129,-0.0011207728113718,0.00292952533582591,0.00103055052736845,0.00418760461997314,0.00663567772410345
"2615",0.00221291182254579,-0.00153566618239243,0.00132028854696165,0.000971350902358781,-0.00672771078098811,-0.00261878742548882,0.00228619303970068,-0.00205841951537411,-0.00633864042804599,-0.00329593395865624
"2616",0.00233270404097508,0.00153802808010273,-0.00150686300614977,0.00388065529372561,0.00563062907524992,0.00206301987351432,0.0067157307698158,0.00386673419670092,0.00394495554763252,-0.00198416790706935
"2617",0.00477948742797962,-0.000877513062653712,0.00264103499499724,0.00483202145606354,0.000324564349726941,0.000561485251247662,0.00213950613009928,0.000256917626584974,-0.0010868489165885,-0.0218687617841493
"2618",-0.000206668016092593,-0.00483096417923123,0.000564488212755565,0.00360670032941268,0.0017036278014988,0.000654391883456729,-0.00615426242030892,0.00154036514386147,0.00887176074141882,0.00745254240077342
"2619",-0.000868846887829511,-0.00154447624247656,0.0020684624714169,-0.00527081863321344,0.00494001350666329,0.00252360430586362,-0.00391764665694505,0,-0.00331841709541714,-0.00806996786866232
"2620",-0.000248401954317523,0.00309380450396968,0,-0.00770702315440031,0.00249822309274905,0.00046600674511188,0.000253755661238309,0.00307648782469361,0.003995372099179,-0.0108473798076169
"2621",0.00795214927057897,0.00638912189402641,0.00900714540388581,0.00849504035005322,0.000104935024794361,-0.000522497807118216,0.004058759444451,0.0091998899241359,0.000829033307186977,-0.00685405688185781
"2622",0.00332858610473541,0.00656751302272185,0.0210154441917105,0.00505429932250734,0.0118404029696078,0.00438837532835312,0.00985350826187226,0.00734359685123498,0.00737243201315074,-0.0048309230214546
"2623",-0.000737188870168159,-0.00587216209185215,-0.00382511337423874,-0.00119745222664014,-0.00620924147308533,-0.00167327916717031,-0.00312722246091557,-0.00276511091416909,0.000986777395059812,-0.00554777457712019
"2624",-0.00319692098143554,-0.00371912204573244,0.000731457324525175,0.000479555135020293,0.00544679362837686,0.00316604085498073,-0.00501964947430056,-0.0015124381856203,0.0112543741578648,0.00697340510093514
"2625",0.00185030868788827,-0.000219674862131591,-0.000365461342886508,-0.00119802594028151,-0.00477996806074932,-0.00185640245590724,0.00416212165033691,0.00403925731194343,-0.00528026816052429,-0.0138503695092584
"2626",0.000492395389298572,-0.00373363011934547,-0.00237609515013826,0.00599783752094352,-0.00264174617448731,-0.00158118261733431,-0.00163295243084316,-0.00402300735008854,-0.0065332382164125,0
"2627",-0.00151758678810088,-0.00286614799435791,-0.00897755287466784,-0.00763166247884495,-0.00152508020756958,-0.000931330654719842,0.00641594532922718,-0.00732143992050971,-0.00912454567818255,0.00561797306157019
"2628",-0.000205668382216362,-0.00508505897129208,0.00314274417266014,-0.00528718128341021,-0.000321302041646931,-0.000186421852407248,0.00662507031609594,0.000254311695897513,-0.00149328022653661,-0.0090782320655145
"2629",0.00489005689783606,0.00577768492275066,0.00552897364170146,0.00483202145606354,0.000160733124823897,0.000372843539189871,0.00211113638022731,0.00991606467621819,0.000997025581613187,0.00422841721504996
"2630",-0.00126764049651074,-0.00176755775347281,-0.000549822144217837,-0.000240469395841658,0.0154365174549247,0.00521994391529002,0.00322165111829698,0.00251790216787939,-0.00547811241339369,-0.0175439077995795
"2631",-0.00192439925198606,-0.00996012052693007,-0.00971954406548459,-0.0103415704258528,-0.00158331106407483,-0.00176161148149201,0.00345867477939499,-0.00502300476757667,-0.00417292605575026,0.00428580271427803
"2632",0.000218532752400913,0.0111781638296309,0.00407414494931224,0.00170112571676539,0.00198230314850489,0.000557239361428818,-0.000615561289197819,0.00349131064587405,0.000167582970164393,0.00426729339038379
"2633",0.00832503562759501,0.0037587883798893,0.00313542515924392,0.00994660784732915,-0.00142467144116298,-0.0027853488121079,0.00172417372603184,-0.00126985101630639,-0.00762523906905432,-0.00637392368741607
"2634",-0.00674417991786769,-0.0104541738453655,0.000333070577655414,-0.0110526659652341,0.00895651128249186,0.00251362793350896,-0.00331982528865304,-0.0162723550814567,-0.00211095161698893,-0.00997862781066583
"2635",-0.000246865094231441,0.000226745139454865,-0.00147981428040611,0.00219626176016274,0.0020423951848898,-0.0000925896100418822,-0.00394737926637834,-0.00258496419557419,0.00287694195295307,-0.010799137029343
"2636",-0.000452793039619315,-0.000906651047564044,0.00203778215706785,0.00511305472846058,0.00219499264210965,0.000928877079207968,0.00198140639612721,-0.00414584276525587,0.00337496633584977,0.00145565913800816
"2637",0.00119445063776991,0.00340289656949011,-0.000739467461176035,0.0053295160771758,-0.000469140903557541,0.000278269798414277,0.00395540957677776,0.004423537632122,0.00428861426654237,0.00436033063266361
"2638",0.000657965717646203,0.00339133141627124,-0.00277521627620314,0.00963861707007663,0.00375599024889328,0.000834735609733572,0.00640246945553025,-0.00207260097979423,-0.00895921460269622,0.00217088652750053
"2639",-0.00805614706770452,0.00247855429351662,-0.0024119906787734,-0.011694509905794,-0.0106814397037743,-0.004912460346294,-0.00591202321381235,-0.00519231055488978,0.00380193474314017,0.0115524115461247
"2640",0.00895027906706436,0.00741745077467382,0.00446340623746888,0.00772763621685946,-0.00330968297342948,-0.000931330654719842,0.0013654757993431,0.00104401347255623,0.000757545673891968,0.00642396808240298
"2641",-0.00878886721284577,-0.0111556374087673,-0.00999796049397828,-0.0127004867187803,-0.00838142819163823,-0.00372930296919149,-0.0109113002869501,-0.00469220913040413,-0.00487806551929248,0.00425518775965816
"2642",0.00186450581643038,0,0.00336629655935172,0.00461156198440893,-0.0023124507067156,-0.00233966533470698,0,-0.00209536914389596,-0.00253552231237308,0.0204803110442378
"2643",0.00169572252073258,0.000451144134383741,-0.0048462045988884,0.00579850714410979,-0.00321958028132907,-0.00367274195660161,0.010655923150221,-0.00892408081069085,-0.0163531693701027,0.0103806233302839
"2644",0.00231199121075032,0,0.000187325291417073,-0.00192171882020531,0.000240804198520905,0.000754235821156968,-0.0112875592058931,-0.00158875351704613,0.00370403148260934,-0.015068498558463
"2645",-0.00914443634169615,-0.00360851187055511,-0.00730348726334618,-0.0120338357064251,-0.00827364240109307,-0.0018843944162148,-0.0174382827773484,-0.00503986300930548,-0.000429076564428699,0.000695472358283933
"2646",0.00648511644382244,0.00203712659381439,-0.000565924720095867,0.0019489770228871,-0.00599372184211855,-0.00160459322848761,0.00485173071115463,-0.00106658976957175,-0.0102172404033893,-0.00972898790088284
"2647",0.00107382520009258,0.00225896019470495,-0.00264249076257728,0.00948207253055777,0.00146674583899586,0.0013232872975637,-0.00736978205259475,0.00186815765733783,0.00164817836266629,0.00421046853524154
"2648",-0.000742625766428251,0.00135227692297391,0.00681312513095378,0.00818880645419928,0.00170866062530717,0.00132209209489242,-0.0011517957465188,-0.0061266042863749,0.00129905602061964,0.00978337842656662
"2649",0.00751487594901779,0.0085527808607917,0.00695485603107082,0.0193502470111708,0.006904548005634,0.00292319498838478,0.0125594133671127,0.00696861741539623,0.00354606460267948,-0.00484429563586741
"2650",0.00168009703413263,0.00424005236829084,-0.00130681187298121,0.00492153332945788,-0.00629264680952679,-0.00103448872020129,0.000379460445425028,0.00452505051216945,-0.00180986815314899,-0.000695400785539535
"2651",0.00466420456398176,0.00622222865798649,0.00243002459522756,0.0125932950498795,0.00121789206989686,0.00141199866480202,0.0101213825590594,0.0135132387643344,0.00820235710585404,0.0111342268915033
"2652",-0.00012234653155585,-0.00154596213071279,-0.00130534983269148,-0.00460612645194536,0.00275689953960367,0.00122175824304849,0.00400821963546361,-0.00235275774854049,0.00445323296531375,-0.00344110942841314
"2653",0.000529629802261455,-0.000884792033848725,0.0052279084352771,0.00300780655435351,0.00873281068962539,0.00366115233709641,-0.00249506108216058,0.00943385247189577,0.00699121828807892,0.00414366093869045
"2654",0.00541395155582158,0.00199245429671646,0.00408614230806226,0.00830448083314583,0.000401010737938634,0,0.0080038748606559,0.00700935821029058,-0.000253992039166984,0.00894087224434292
"2655",0.000445382367051383,0.00552375081196099,0.00369958455073349,-0.00114389165405271,0.00288453916045928,0.000280532295924063,-0.00397011905296651,0.00438263882764089,0.00135497965184661,-0.00136337802319941
"2656",-0.000890303325772779,-0.00593263408804556,0.00184300323888786,-0.000687165702332515,0.00423457198991639,0.0017765119146691,0.00211735769348032,-0.000256800260155288,0.00862655630288489,-0.0136518315761254
"2657",-0.000243129437243139,-0.00309475422773042,-0.00202359548439546,0.00297961647388267,-0.00389851642649652,-0.000653347382286951,-0.00261008638566529,0.000256866223468322,0.000419218507140329,0.00207609617564697
"2658",0.00243089007858321,0.00221721749713111,-0.0035022718804858,-0.00251370112610649,-0.0130193616527452,-0.00560399070970541,0.00124623795434942,-0.00154009488397822,-0.00326879562934856,0.0110497861959944
"2659",0.0000405202186370968,0.00774349223009407,0.00332965540549091,0.00824743036566788,0.00161861734055058,0.00319360216291553,0.00535213501559229,0.00437021493744671,0.00807264561171617,0.00956278073642225
"2660",-0.000929703581005858,-0.00461039478188519,0.00331858611739921,-0.00545331110682934,-0.0049284615472579,-0.0015915231553949,0.000866757505772142,0.00179171353858809,-0.000750717402837386,0.0060892964033703
"2661",-0.00117291672223863,0.0011028249333056,0.00294006932272239,-0.00045695917852806,0.00592708013799181,0.00168786307466329,-0.00210288434061268,0.00383242325680166,0.00751315629423854,0.005379955507687
"2662",-0.000567078736324,0.00264375331893341,0.00329783602130762,0.00114292021420259,0.00121104329160149,0.000280485563450839,-0.000123888665608196,0.00152682426159512,0.000497124857119502,0.00602005367344782
"2663",0.00222877156142887,0.00483409691040482,0.0058437650064993,0.00296797726595432,0.00702084201118258,0.00248420552466944,0.00446307294267911,0.00330379597043007,-0.000828140786749532,-0.011303174426881
"2664",0.000485324690663091,0.0010932522901228,-0.000544752151579231,0.000910392216531886,0.000561702186401947,-0.000935249541174965,-0.00629487235252124,-0.00253278438853488,-0.0020721093730276,0.00201745736003356
"2665",-0.00193983462242653,0.00152917311474354,0.00254312737930085,-0.00409360607134579,0.010344046176928,0.00346301223782874,-0.00347769770983575,0.00126948624761236,0.00157802322960099,-0.0073824498756202
"2666",0.00182201684082361,0.0019629041003657,-0.000906002299686959,0.00365397929017908,-0.00849235468273291,-0.00270461856843585,0.00336548966033057,-0.00202897309091632,-0.00779495838112476,0.00202830017005384
"2667",0.00185916021284704,0.00108842145095078,-0.000362626104956965,0.00682582081309713,0.00112106430495018,0.000560812698353175,0.000745193979066361,-0.00355795986248686,-0.00117007937868652,0.00202433339157682
"2668",-0.00246091004639193,-0.00652321450850202,-0.00108852208462795,0.000225927633690004,-0.00359808857486654,-0.000840792311486038,-0.00546178541736997,-0.00382533868860191,0.00292861680313594,0.000673322171594659
"2669",-0.0000405464368633535,-0.00131318531813907,-0.00617505821641651,-0.00903739219642774,0.00545625603421018,0.00121605732111418,-0.00174736876171666,0,0.0120974218913947,0.00672959153000807
"2670",-0.0141151870992114,-0.0149024642584514,-0.0104166477646286,-0.0237118314156815,0.00853967143578038,0.00373698816478552,-0.0076269032898072,-0.00972852474530506,0.00741901751576979,-0.015374396255745
"2671",0.00147684350926847,-0.00200220586330568,-0.00147743278336276,0.00233513146342279,0.00047480204979089,0.00111723757288695,-0.00478765909745016,0,0.00474594554247565,0.00339445675241579
"2672",0.00991303901511231,0.00735607690976225,0.00739787920455792,0.0102519458593544,-0.00514094935399367,-0.00241749503769084,0.015318362448536,0.0067216116864699,-0.00708529190418361,-0.00879568904694039
"2673",-0.000121470223129028,-0.00110638888410386,-0.00128514204825214,0.00115312497568842,-0.00421378278292639,-0.00298273083623413,-0.00286798231787422,-0.00487891477338764,-0.00770993286925747,-0.00477816212774163
"2674",0.00174420290608479,0.0053168636837988,0.00330884513881236,0.0103662212629232,0.00367250971281785,0.001869761447437,0.00437681949453972,0.00851585398150445,0.00735658768333813,-0.00274344684758798
"2675",-0.0155907969304365,-0.0125605535390149,-0.00677902923264029,-0.0127679092238284,0.00747765338958151,0.00354586608231688,-0.00684785136547017,-0.00639713899049277,0.0050873470479853,0.00275099405355195
"2676",-0.001563063951313,0.00066941389222186,0.00442717827596106,0.00854485447402453,-0.000236773994166328,0.000185958873014647,-0.00739610122696432,0.0038631434876979,-0.0015511062380783,0.0178326868731391
"2677",0.000782689445435247,0.000892166086847945,-0.00220387117901344,0.00366389608855489,0.00244819763683846,0.000650779570066984,0.00896711059857647,-0.000256545660889618,0.0037612345765845,-0.0121294223954782
"2678",0.0104569848566343,0.00579308215839802,0.00202465469229773,0.0111797544642687,-0.00386048458467136,-0.00195121731274206,-0.000876416936580138,0.00179618830258299,-0.00448031110328595,0.00272854600406491
"2679",-0.00358537342453069,-0.000221474425783241,0.000367502231693129,0.0047382343806861,0.00680173633103909,0.00344430562773379,0.00826854054181525,-0.00076857684043663,0.00376400461307602,0.00884355670473025
"2680",-0.00233056848417945,-0.00132948009086731,-0.00514143424741553,0.00314387754510492,-0.00369205976041032,-0.00157711805359073,-0.000993950543650701,-0.00358847897656034,-0.00309771750383503,-0.00067436901525264
"2681",0.0023360127218075,0.00710008065417589,0.00332226120894186,0.0058203937560577,0.00386339238071387,0.00167225757066247,0.00472642237856191,-0.00128638896933564,0.00367975301594758,-0.00202419449601332
"2682",0.0000409940798764552,0.000220447264182466,0.00110375992307388,-0.00356097789903687,-0.000628371061380029,0.000927710253414205,-0.00507555636010293,0.00309083528100529,0.0158872741712119,0.000676053664256049
"2683",0.00114480798367689,-0.0039649365739709,-0.00202136438339917,-0.00178703359473431,0.00322218615684178,0.00231671669110223,-0.00149313356401382,-0.00205428961222842,-0.0021654021627171,0
"2684",0.00473751152334656,-0.00176916853720899,-0.000552456142521085,0.0015663596517288,-0.000313149527788936,-0.00083191355853196,0.00535836116427468,-0.00154393501013506,-0.000482213478254612,-0.00743240066882345
"2685",0.00601615564896374,0.00731073903429103,0.00792194207127794,0.00156400693725933,0.00297758004009374,0.00157287243067605,0.00644495358563435,0.0108247815007008,0.0117401012243479,0.0279101820157066
"2686",0.0014142708855589,0.00219917529664015,-0.00402118398679541,0.00736118488546933,-0.00764879695619192,-0.00294253048614712,0.000123287058183097,-0.00382460609005097,0.00190747099030353,0.00132448516535044
"2687",-0.0071821404264969,-0.00636385597940403,-0.00440448726028564,-0.0130648260906563,0.0158576670878843,0.00696017901846724,-0.00209320696574045,-0.0010236043299422,0.0111058307330769,0.00198403176737982
"2688",0.00341368787132268,0.00706705538908059,0.00423969475771035,0.00650671054946694,-0.00613539637621929,-0.00239610583733818,0.00197406723667282,0.00614899246527667,-0.00509964698807197,0.00990112731437764
"2689",-0.000121487816056365,0.00899134422955505,0.00587372084763427,0.00735606894607921,0.0102369065728709,0.0043418006429099,0.00652727280430021,0.00814865284864807,0.01040932908145,-0.000653653071059468
"2690",-0.00117475283426083,0.000217381613279555,0.00310216808845687,-0.00663854794853813,-0.00216573621183647,-0.00073593175786435,-0.000611807070292736,0.000505215887647514,-0.00124876292637321,-0.0111183607233376
"2691",0.0106659291104247,0.00760530121004033,0.00454798718149863,0.0133660913594706,-0.0119382906303342,-0.00570698437950201,0.00844762328420368,-0.000252707043361333,-0.0139095021183909,0.00198403176737982
"2692",0.00337086527234964,0.00452867700361281,0.000724239609146249,-0.00109910788567935,-0.00525629731147859,-0.00240705417005271,-0.0100763880123922,-0.00429287365259745,0.00293205479147218,0.00264029608816352
"2693",0.000479705498636296,-0.00601114707146733,-0.00199048514876032,-0.00528169467953077,-0.00394355055891771,-0.00204122844166521,-0.00367910712319353,-0.0073546138152264,-0.00750629752696419,0.00460829992672163
"2694",-0.000319628975010366,0.00323999414752785,0.000181270567237268,0.00265477356266919,0.00411748699419245,0.000185618766328943,0.00615437788310813,0.00204391421407935,0.00437865612309007,0.000655366512221311
"2695",0.00134605348910899,0.000430433024755539,0.00145030386808487,0.00595758046852568,0.000394257243778062,0.001208970728799,0.00415958475025913,0.00324024336909634,-0.0049936983197939,0.00458415661069123
"2696",0.00212703050524565,0.00193673872284594,0.00018105173503602,0.00350961648955161,-0.00575445035913369,-0.00390042989203254,-0.00536075078606413,-0.00281964803228241,-0.00932046530168462,-0.00130376311982083
"2697",0.00100100912744261,0.00472508066552235,0.00579178464142815,0.00218574697991358,-0.00245787038877632,-0.00111844812783557,-0.00771665895505869,-0.00308481050558718,0.00209072047209125,-0.00195826488688433
"2698",0.000360029797722428,-0.00299268826108634,0.000360029187075783,-0.00458019265334353,0.000715385602792828,-0.00195993451458776,-0.00246899256314503,-0.00257884422901922,-0.00802439396506838,0.00850230752397341
"2699",-0.00267932995996034,0.000857570146966413,-0.00395766060387204,0,-0.000555808190463636,-0.00130900674272483,-0.00321735593427896,-0.00698014871686758,-0.00760397166468274,-0.00389106408858941
"2700",0.000200532404304621,0.00214226403897899,0.00108362642400173,-0.00569669175553689,0.00286062531972386,0.00177899474099985,-0.00595896587875766,0.00442577488138074,0.0045647049233779,0.0039062636106455
"2701",-0.00204465135117038,-0.00769564102362152,0.00216496406851419,-0.0169678076065254,0.00626012689525202,0.00299078994157131,0.0053705189091291,-0.00544304218010849,0.0104673890046638,0.0168611887231829
"2702",0.00060264486762418,-0.003015897525809,0,-0.00268988508625156,-0.00181135477920735,-0.000838387142237385,0.000275374474416168,-0.00208497785656325,-0.0111619690930858,-0.00892858080554015
"2703",0.00389436280798905,0.00172848199847153,0.00198018871901695,-0.0035964630822034,-0.0150677976929461,-0.00512996433993695,-0.00801605752552281,-0.00443989301806158,-0.00942013975491429,-0.00386108364400783
"2704",0.00119969117988838,0.00345135275755637,0.00071874218750767,-0.000676804452399815,-0.00296344820312155,-0.000187361867199365,0.00744958521817973,-0.000262358724170242,0.00188552217038396,0
"2705",0.00351512393464914,0.00752367715249536,0.000179499598359056,0.0115125621346592,0.00224916994671709,-0.0012191366214851,0.00112790979729338,0.00708467255114398,-0.005155036454914,-0.00516788856168493
"2706",0.00433864339840495,-0.00192021011229326,0,0.000223176777647716,-0.00183121944058351,-0.00113758692991606,-0.00200284741290913,-0.00234476912830739,-0.00666232099584918,-0.00844151018349193
"2707",0.00214011869196429,0.00320649177392851,0.00592340965352123,0.0158409266284434,0.00096566881407556,0.00141230140735016,0.000752493193792336,0.00470080794361638,0.000496853535568054,0.000654869887072751
"2708",0.00118648536200894,-0.00170463500204854,0.000178467133575166,-0.000219552268222012,0.0000803357890986067,-0.000282169646196206,0.00639274049793248,-0.00519888074226238,0.00281383757653186,0.00130894998339981
"2709",0.00592508566819205,-0.00128067097656459,-0.000535098558641312,0.00746929959765419,-0.00377792974110458,-0.00103414582849981,0.00311361592911119,-0.00130659011641931,-0.0053643724579413,0.0111110931727056
"2710",-0.0011388625161648,-0.000854914409601504,-0.00053559246097612,-0.00501523323257624,-0.00282386071648533,-0.00122372718809649,-0.00360072214469997,-0.00183114735350287,0.00472949729661876,-0.0155139513659167
"2711",-0.0016510961641335,-0.000427858036726847,0.00125030997393893,-0.000657427157144674,0.00315556734609346,0.00113070065622356,0.0019938345126076,0.000261903496820759,0.00817578687507758,0.000656522276818006
"2712",0.00263835075994856,0.0106997660220938,0.00713511975942738,0.00986846565207644,0.0016131981152081,0.000376527809505811,0.00136767520928371,0.00707548306739159,0.00262123193608743,0.0118111334310549
"2713",0.00157098553505208,0.00254073425080903,0.0051363164192284,0.00456020562203552,0.00193263341694938,0.00112915826902782,0.00422294574909854,0.00572452952935776,0.00318626628780616,0.00194549867153038
"2714",-0.00149009263045885,-0.00190072145999209,-0.0012335099777796,-0.000432456584116392,0.00425987424791585,0.000940088429009611,0.00655443471634887,0.000517614316628112,0.00081438227205477,-0.00129448070386373
"2715",0.001217435171601,0.00169282474253052,0.0123500917613661,0.0090831481860445,0.00720288071920838,0.00338000787704651,0.00221126885882539,0.00284468469636345,0.00756775170939661,0.00972125587305173
"2716",0.00133366365248699,-0.00253485351409566,0.00453119444127137,-0.000642821737533272,-0.00071526328981697,-0.00168428116327779,-0.00502600119130103,-0.00128931500312801,-0.00686479567113552,0.0025674912770961
"2717",0.000704987502999632,-0.00381209348814171,-0.00104095058667075,-0.00514709135466074,0.00127216397329533,-0.000375044373884803,0.000862485105386002,-0.00103275294311445,-0.00683096684694662,-0.00128045807361343
"2718",0.000978541346826844,0.0042518317944904,-0.0010419619124461,0.00237119135542763,-0.00659138202931719,-0.00253181271792269,-0.00110802417046207,0.00439374532233971,-0.00376647024727261,-0.000641082861988718
"2719",0.000273782593481764,-0.00169344878563726,-0.00226011949819427,-0.00881717815589933,0.00175878875305968,0.00103420824150913,-0.000739420008804004,-0.0012867524841671,0.00591765440811454,-0.00448993064839287
"2720",0.00516055117125624,-0.00296866680820851,0.00226523920949973,0.00368849810534222,-0.010613708996479,-0.00413223016953457,-0.00320685321403091,-0.0043801609575671,-0.00637305340610395,0.0051545684159735
"2721",-0.00388957865986517,-0.00319010198978931,0.0024337926118243,-0.0079983600225918,0.00177460452744382,0.00094305963835728,-0.00470168700452067,-0.00879923091807633,0.00156238794866881,0
"2722",0.0017571125734348,-0.000640085588587191,0.0083247535055162,0,-0.00619961170291117,-0.00301519950884999,-0.00497290220713131,0.00156659935921799,-0.00385879300840419,0.0102564681117521
"2723",-0.00494994464582943,-0.00106741479535877,-0.00808393052228928,-0.00217891345665189,-0.00478030445497191,-0.00160619096103531,-0.00387293816677581,-0.00782062106895687,0.000164806722742883,0.00126895282363715
"2724",0.00129255204497492,-0.00235098541813294,0.00537537664709609,-0.00677024384347402,-0.0033376159745051,-0.00132524158190916,-0.0061455135092563,-0.00157644681933555,-0.00840540598937634,0.00443606490635928
"2725",0.0081761334472632,-0.00171376438782134,0.00758882487610313,0.0145117924904039,0.00661601883951346,0.00322235265184356,0.00454317787061553,0.00447362056416933,0.00473697324462785,0.00504724945748625
"2726",-0.00372492780295541,0.00579398387426822,-0.000342392944072789,-0.00628511990967673,0.00957482791219455,0.00359005787312672,0.00213544325787307,0.00104815353069121,0.00190235728862942,0.00251101593966951
"2727",0.00155769570660635,0.00512059140176113,0.00428092551990877,0.0093783342605962,0.000321412346220962,-0.000658768319409142,0.00188054860239961,0.00680426478035256,-0.00379756469406989,0.00250479097826695
"2728",0.00132219191087768,-0.000849084087615082,0.00562655395007772,0.00518590119045514,0.00445247626068923,0.000603605978459987,0.000750610102697724,-0.00441899618615471,0.00364633303466189,0.000624536740310377
"2729",0.000388510252994578,0.00254927756648526,0.0011868716510488,0.00128986236867057,0.00440901833956064,0.00132006732700995,0.00625148075369242,0.00391626599708772,0.000660564770369465,0.0062422403245177
"2730",0.00333861698691029,-0.00254279527553314,0.00237078620390263,-0.00515243049307967,0.00271366067523626,0.0016004750933738,-0.000621001953927336,0.00130038100577012,-0.00470335003377598,0.00620332494232834
"2731",0.00154763907309974,0.00212449088254441,-0.000168826621252616,0.0112213935661305,0.00374050891783195,0.00122266006481309,0.011562789512126,0.000260108352175381,0.00853920555780463,0.0191123283471131
"2732",-0.000695357512788486,-0.00826800488720703,0.00794188499120119,-0.00640196184770436,0.00420286194731245,0.000375107752076831,0.00712864462946272,-0.00259680144991647,-0.00361695842799903,-0.00604964843524292
"2733",0.00170090538944323,0.00064120019401237,0.00620282214958023,0.00472488009993577,-0.0022109779776992,-0.00121980412227918,0.00671228965696713,0.0093723981910796,0.00346504416685955,-0.00182590324516907
"2734",-0.00362760686573627,-0.00704954671308577,-0.00833056360075968,-0.00619903968062896,-0.00284886873098233,-0.000376331122240336,-0.000363659495808744,-0.00232142717752781,0.00411082802213669,0.00182924326638534
"2735",-0.000310142678561887,-0.00150614305484587,-0.0073925447997174,-0.00430212064835933,-0.0150795559430835,-0.00507661559159767,0.000606400496201198,-0.00180949318266743,-0.00818799659841141,-0.00182590324516907
"2736",0.000930020570554912,-0.00452486790355899,-0.00440074004351609,-0.00216027241823902,0.00209525230337371,-0.000472261362645221,0.00363587481043615,-0.0049211226106739,0.00148601506198331,-0.00304873877730882
"2737",-0.00232253923801684,0.00216435556430206,-0.00527037140159448,-0.00671142736248043,0.00675454906963058,0.0014181546309191,-0.00156992925108157,0.000780652350691247,0.0020608359090073,-0.0134557875869372
"2738",-0.00500526721305727,-0.00453552425106352,-0.00734920417788165,-0.00523111335944226,0.0108625925717469,0.00358722526520405,-0.00858734102588832,-0.00130013407844909,-0.00123390920095268,-0.00123984494504614
"2739",0.00850093150441289,0.00650913280212673,0.015495915228789,0.0208151314156375,-0.00869153354737928,-0.00253969485989181,0.00670992797304915,0.00937474647342129,-0.0000823820086522931,-0.00310368377575998
"2740",-0.00293869721528961,-0.00129346416202558,-0.00491691432785057,0.00493658169677902,0.00741260462004156,0.00132000643502028,-0.00460492093383147,-0.000257781793636336,0.0120263507079679,0.0161893255167598
"2741",0.00170631451932213,0,0.00494120983327684,0.0051261126525759,-0.000395612699329639,-0.00160108623284372,-0.00206981533016792,0.00258047337375955,-0.0126160099901025,-0.0079657033931777
"2742",0.00654276087193195,0.00539589490704517,0.00915568792330301,0.013387028465373,0.00316615416543242,0.000188715715695453,0.00719793752125075,0.00592028633606212,0.0016487017005804,0.0067942881877463
"2743",-0.000884411679163755,0.00364977338403438,0.000672059207656561,0.00251641276956938,0.00323510080911915,0.00320655259777292,-0.00278590723573247,0.00230276962497822,0.00921730706580015,0.00552146022906941
"2744",0.00230956493616397,0.00919783692563358,0.00822698330490157,-0.00209156922889275,-0.00275273573563362,-0.000845888444582887,0.00206494428240123,0.00459547319545628,-0.00252790514216528,0.00305072465542766
"2745",-0.000499115009775841,-0.00635868282490559,-0.00432970643716102,-0.0146720351692161,-0.00141964776657533,0.000658667393373058,-0.00412148588644468,-0.00101648109042951,0.00416940810987576,-0.0018248551037251
"2746",0.0101447564382307,0.00639937441710181,0.0030105387051973,0.00744538152339858,0.00134258398644782,0.00018781347762542,-0.00219065359896964,0.00432468941900233,-0.000162859233691082,-0.004265696046719
"2747",-0.000608636966939469,-0.00402713102891006,-0.00200094299621689,-0.0158362644035293,-0.00985879391358091,-0.00319630348253774,-0.00121990199936295,-0.00658553559365116,-0.00626982340639715,-0.00673198010526599
"2748",0.00875503200760042,0.00106393763301682,0.00100231855219102,-0.0109419960183423,-0.00334546234619393,-0.00311246235815843,0.00109913337101863,0.00484437140640726,-0.00770241717713527,-0.00431300522668032
"2749",-0.00207546745955212,-0.00361380368276387,-0.00450665765982816,-0.00563975450480392,0.0134945274166243,0.00369567112105518,0.00183017134890329,0,0.00404622632611429,0.00866337563776698
"2750",-0.00121007184978739,-0.001493610795818,-0.0105632806845122,0.00196338804343843,0.000474234934866313,-0.000471870174931666,-0.00767200087346809,-0.00380608318027376,-0.00337195504143284,-0.0122698975885782
"2751",-0.00359654397470033,-0.00363233592188728,0.00254175245177413,-0.000653203850350836,0.00497576796373789,0.000755364692971217,-0.00589015929669023,0.00382062479604817,-0.00709688067337855,0
"2752",0.000190017772597306,-0.00171569571069508,-0.00371864028795643,-0.0135076610327362,0.00345790871189577,0.0020760743846433,-0.000370193600061519,0.00177621631805036,-0.00207779255319152,-0.0167702126206949
"2753",0.00315295753483347,0.00257794308514225,0.00644717482270107,0.00287087171309008,-0.00783181852900683,-0.00178953087919909,0.00407521543719214,0.000759572353670634,-0.0131590072457732,0.00315851657128929
"2754",0.00545325091889426,0.00514246477913072,0.00472020466519107,0.0116715104086151,0.0000786893519102438,-0.00075465099953953,0.00332048726733647,0.00379678147675255,-0.000084353111390878,0.0050378444325565
"2755",0.00301291346610477,0.00191864266164332,0.00335582109086285,0.00500659436553619,-0.00205215944933568,-0.000660807074430392,0.00110306616685074,-0.00176490012569663,-0.00396692258692799,0.00250629588749507
"2756",0.00176473717895553,0.000425419325789322,0.00183926174033688,-0.00671433479056294,-0.00039545954160336,-0.000850436486029116,0.00404058196558688,0.00303095653149876,0.00118634012056029,-0.00875007309041997
"2757",-0.000112305910477173,0.00212677341372558,0.00400608836143057,0.0119931403032116,0.00751721992611176,0.00406613810886136,0.00207345796979563,0.0095696085028385,0.0086330595237738,-0.00441362391405054
"2758",-0.00408615374030363,-0.00594228116818696,-0.00465521166382354,-0.00732608368912335,0.00424084273820791,-0.000376645282451293,-0.000608527017794902,0.000249229701419162,-0.00201391293134034,0.003166583158283
"2759",0.00832734882031683,-0.00106741479535877,0.000501291948905802,0.00217058841630391,0.00375385377517512,-0.000188209206987477,0.00414013803120916,-0.000727081656357709,0.00210207685192976,0
"2760",0.00634129483681778,0.0132506709665603,0.0120198822829269,0.0112626884435656,-0.00911564560566225,-0.00226149766946193,0.00557846418342467,0.00978431572030947,0.00461489343849641,0.00441919659547785
"2761",-0.00384048295960437,-0.00105458147505533,-0.0101458396159084,-0.00528339545669521,-0.0129740440092477,-0.00453383677124519,-0.0192564878845153,-0.00322971950847373,0.000751666230226267,0.00754251726589228
"2762",-0.00052391134091534,-0.00401184797514831,0.00134200465776813,0.00131139960355808,-0.0110728630721426,-0.00294094145477231,-0.0104387934472975,-0.00174504740838666,0.00267066432982821,0.0056144599261303
"2763",0.00205968961940384,0.00420360710696288,0.000670094257276821,0.00654880694077398,0.00582828268786417,0.000705273608409884,-0.00364179319937208,0.000749450115848482,0.00141500750303813,0.000620211184653829
"2764",-0.000261585885439342,0.000850016918630292,0.00468778225086552,0.00845803333930872,0.0013644499042611,0.000380756385184089,0.0063019680507086,-0.000499200331025018,0.00523650578067514,0.00433987205688369
"2765",-0.00119634758737253,0,0.000499890769661393,-0.000860218997046358,0.00296540068842566,0.000380913138490646,0.0048850010423136,0.00149784798730468,0.00686286577041728,0.0148148021084444
"2766",0.000486602554070181,0.00148614518196144,-0.00133239348787073,0.00258290183013665,0.0130255353901658,0.00428215342332838,0.0036142419516807,0.00648069247049876,0.00377766289999992,0.00243299406141095
"2767",0.00205751465247217,0.0023319515052278,-0.00233485635438169,0.00687002427882644,-0.000867965457523323,-0.0012318894672344,0.005837103373036,0.00346692055979458,0.00507236345236772,0.00485430284159838
"2768",-0.0037705680264718,-0.000422858558315142,0.00183884217638464,0.00469072704196005,0.00157915453342317,0.0016131713963341,0.000247108243740746,-0.000740436398890876,0.0065120391780551,0.00301940706457482
"2769",0.00715722399981922,0.00677112729687579,0.00600697667984695,0.0188879576339418,-0.0107992308017085,-0.00331542647979477,-0.00506107476522943,0.0059273264347337,0.0121310147653697,0.00481637198410567
"2770",0.00632502386726275,0.00273214007647793,0.0137667762280753,0.00958139168865246,0.0047811135111977,0.00104542806093511,-0.00161291129984953,0.00564692826249846,-0.00263685173572759,0.00599165342118746
"2771",0.00421490324968188,0.0121568360944448,0.012270838604596,0.00495151648830894,-0.00015855992588687,-0.000474579796318264,-0.0156581833398922,-0.00146470578995284,0.0051273754206056,-0.00119116894609306
"2772",0.00666425047274832,0.00683364222450678,0.00274784297887964,0.00862244315219929,-0.0028556653606856,-0.0012345836317692,0.00101020080183711,0.00440093813557363,-0.00103616292871167,-0.00357789130999808
"2773",0.00182851142473517,-0.00267369888629687,0.00580272828007611,0,-0.000636470974227921,-0.000476014846736983,0.00567525841622496,0.00024323687121508,-0.000159610625395157,-0.000598312713800175
"2774",0.00226340551641635,0.00144354361665844,0.000640941923124361,-0.00162827505471785,-0.013372449504117,-0.00475726982411573,-0.0115374313177724,0.00146021556165055,-0.00462848144008432,0.00658673582176394
"2775",-0.00152983001521456,-0.00329497343475904,0.00640628855164738,-0.00632022389305242,-0.00121004948108328,-0.000286512983699416,-0.0121797945117348,-0.00680409737667242,0.00240516309456029,0.00356925525226215
"2776",0.00729607594653392,0.00702487304939758,0.00668356095727241,0.00615510399068975,0.00411973177530722,0.000669452530334791,-0.00346797820440237,-0.00122341539773729,0.00327923700935173,-0.000592638145727076
"2777",0.00651915911587109,0.0133359811795808,0.00316160713810287,0.00958397519763143,0.00168889840736641,-0.000669004663470085,-0.00811915072209568,0.00710420607012918,0.012117322829762,0.00652416725529137
"2778",-0.00341837049285421,-0.00080985092246455,0,-0.00383745901504717,0.00417619120729928,0.000478180378810533,0.00272871792299001,0.00316227042855455,0.0016540564087435,-0.00471419813690632
"2779",0.00953150122026347,0.0044580103220826,0.00803650497152719,0.0131792260399053,-0.00135952058248456,-0.00219851784855285,0.00712685759216214,0.00703219923095966,-0.00809938677517319,0.00118411653188644
"2780",-0.00168055836200265,0.00100859379853291,-0.00844144558312043,0.00120058682051205,-0.00928967541231762,-0.00316146290980024,-0.00977846018292883,-0.00120408638914771,-0.00221973998905778,0
"2781",0.00454946739047601,0.00483682324287993,0.00630616797922201,0.00819500858873745,-0.00525425189756779,-0.00259446467712976,0.00649685628244678,0.00120553796099809,0.00444936433776144,-0.00177407408737407
"2782",0.00813087156112968,0.00681914858436294,0.00422994726844172,0.00574953276824641,0.000975035452622564,-0.000385419229865125,0.00813309990957922,0.00650109431775991,0.0018193640534625,0.00236963602636964
"2783",0.00212285471228202,0.00298791651758346,0.00608418985661019,0.00473092893046201,0.00430277407185331,0.00289177912505489,0.0138300548453236,0.00406721925048203,0.00497431496290068,0.00709240651970733
"2784",-0.000388876275475791,0.00317772580325215,0.000310239713469107,0.008436441647933,-0.00541612101531197,-0.00192229051684267,-0.00353644776639761,0.00619471941448357,0.0121778992157284,0.0105631140112774
"2785",0.000424020878772469,-0.00395955330619924,-0.00480558121648933,-0.000583790104466742,0.00820878514841161,0.00221481903706522,-0.00190144684658655,-0.00331515525623938,-0.00667547144802505,-0.00580700294982217
"2786",0.011577752624262,0.00795067374820091,0.00732095085420004,0.0138213233939251,-0.00370819322424421,-0.00297854396953823,0.000380932865675199,0.00855310771589934,0.000781480028276382,0.00759347409706135
"2787",-0.00662981142890884,-0.00985988468798116,-0.00850468086035794,-0.0151689424511772,-0.0069584206191674,-0.00250557533900275,-0.0128220661588778,-0.0150764929320545,-0.00562199547627107,-0.0028985109481735
"2788",-0.0102570677745681,-0.00677161401397741,-0.0127885779447691,-0.0136478734329019,-0.00586655189711383,-0.00231879118440159,-0.00540130409184403,-0.0047833851380209,-0.00431876724489622,-0.00697676784298473
"2789",0.00049683861911376,-0.000200492232935279,-0.00568722395193888,0.00869728356488575,0.00590117142553548,0.000290755249315211,0.0157744545389751,0.0108145514365519,0.00670346198651117,0.00117094409959151
"2790",-0.00113539092553894,0.00180518407614283,0.00492543728154926,-0.0135214102553071,-0.0144927770581353,-0.00515845205455912,-0.0166750984486523,-0.0116499679460911,0.00329028588656044,0.0099413840415421
"2791",-0.0217697203067921,-0.0248249340158446,-0.0147036564903423,-0.025625622821121,-0.0092792462298108,-0.00370391813706439,-0.0102264610902849,-0.0204474722144211,-0.0131178879376496,-0.0162129851678451
"2792",-0.041822674477441,-0.041264564077257,-0.0473362999805044,-0.0350663270402948,0.00945006025257289,0.00821764786410917,-0.0321737459263193,-0.0351179517259679,0.00253184589391431,-0.00941735710162106
"2793",0.0197025325161451,0.022055608789578,0.0242546535178398,0.032537411960156,-0.00621330882230675,-0.0043666378756777,0.00351353131335097,0.0132348638700877,-0.0104964249901067,-0.0059416896181449
"2794",-0.00542503391076032,-0.0121517417257521,-0.00888003771187662,-0.031512090102757,-0.00950328081521257,-0.00292354075934964,-0.00390536571406197,-0.00979669282439399,-0.00470566289772678,-0.0113568727483593
"2795",-0.0375088918605334,-0.0250263782757043,-0.0296998316249021,-0.0346503930468997,-0.00109400749943345,0.000880121409505774,-0.0294713084084047,-0.0228309091035417,0.00152257391199151,-0.0102780351854992
"2796",0.015021479921971,0.00348042652609704,0.0100890070977537,0.0159771880869231,-0.00631912630711717,-0.00175823153241306,0.0207550400192342,0.00882635476948135,-0.00168031681036196,-0.0146611405460728
"2797",0.0146845000471345,0.0123564729844008,0.0194683948093612,0.0157261160538882,0.00440925042417772,-0.000293181616308869,0.00300207856404078,0.00823507924478606,0.00480889648494576,0.00619967137823907
"2798",0.00248744188125238,-0.00214152809119339,-0.012288319094356,0.00763515035781959,0.00447390756884491,0.00166350082340205,0.00761910189408455,0.00306240770178601,0.00566322870710945,0.00184840363382421
"2799",0.0134960779650217,0.0199570984967505,0.0151311998549366,0.0250473877612567,-0.0110932623774584,-0.0060571649734934,-0.00486069604002293,0.00610725748548169,0.0170526171152821,0.0153751344041695
"2800",0.0127602170027747,0.00736382110611489,0.0048028570492562,0.0205338857239317,0.00339923602970127,0.000294730624811779,0.00990485982908029,0.00354078218768983,0.00116984328690162,0.00181718054121949
"2801",0.000292952969692228,0.00104437526356937,0.0153288818002015,-0.00321937339148226,0.00542066461088586,0.00235839371544877,0.00846419428362455,0.00579614585769561,-0.00327158423151652,0.00181375993405042
"2802",-0.00626126881028621,-0.0110578401470861,-0.00811688823300005,-0.0137262581350066,-0.00438064936269977,-0.00107839063721615,-0.0123900934031869,-0.00501122720061853,-0.0134417084514044,0.00301758450131029
"2803",-0.00497410604521031,-0.00443037781784839,-0.0099835624460114,-0.000818756761560513,-0.0122681989022203,-0.00294391019501394,-0.0165925140718736,-0.00805832788470062,-0.00459437586492994,-0.00120347674362009
"2804",0.00129595493192736,0.00508579802565601,0.00462881484121325,0.000614619998267951,0.00299816309257128,0.00137786866072176,0.00932792519876546,0.00279237838048774,0.00509310026760779,0.00903620732628263
"2805",0.0159394495859047,0.0067467437853963,0.0146454536512883,0.0178096196106146,0.00888182462848053,0.00383336383426469,0.0169885338315083,0.0151898180315773,-0.001266856660328,0.00656719708467035
"2806",0.0116123168324929,0.00649234133248267,0.0129743145991672,0.00925179816444244,0.000338812710309666,0.00117512265100017,0.00347433901927285,0.0107231299533774,0.00245757097239219,0.00533812706251435
"2807",-0.0124866123442812,-0.0158137985185124,-0.0136086758032063,-0.0290953141972925,-0.00143893920557325,-0.00312968320201834,-0.0210412466113121,-0.0217121827869671,-0.0104389089072101,-0.0100296031652974
"2808",-0.0101300623342616,-0.0109935773392216,-0.00876478184338747,-0.01436789291263,0.00635615117146604,0.00235437042262943,-0.00244853891904917,-0.0103403043620608,-0.00103889557353709,-0.0107270933030973
"2809",-0.0145407143088225,-0.010688285261804,-0.0289832271201294,-0.00187402199532738,0.00682645790889236,0.0043032571552033,-0.00313682124063408,-0.0030580862187346,-0.00223999200000002,0.00180720426467462
"2810",0.00515511017813131,0.00108038762708329,0.0112984983392026,0.00417272597268514,-0.008129466530303,-0.0037087496270013,-0.00177839494682441,0.00996927463359421,0.00537201727572145,0
"2811",0.0115577883343745,0.00669111795799782,0.00450235016302125,0.00145445082776519,-0.00270392341617609,-0.00127400238167796,0.011237793994739,0.00202489175458398,-0.00167476674116562,0.00601333289763395
"2812",0.00253512561765912,0.00578908955950297,0.00614198825419332,0.00933604676513489,0.000932002435451995,-0.0000978741296965291,0.00636924919848014,0.000252301787886822,0.0107844623741811,0.00358632258656688
"2813",-0.000366567842238985,0.00255792655055931,-0.00841451897540613,0.00102772638657789,-0.0011004285478643,0,0.0051169745074342,0.00505069551516635,-0.00640162812298772,-0.0107207044128849
"2814",0.00483930743034899,0.00170114136873956,0.00615648886184061,0.000205378129416678,0.00576231672170557,0.00206029921632922,0.00509104221105616,0.00427124564813286,-0.00238627901379029,-0.00602051145286409
"2815",0.0174022378284135,0.00466995777091506,0.00248054437485656,0.0213507719225967,-0.00657176923279246,-0.00215390019209605,0.00626504379953108,0.00150122073314418,0.000956809136609893,0.00969115162118062
"2816",-0.00125525503855684,0.00169015195142141,0.000989859539724192,0.00241211422424925,0.00576692402249823,0.00235440842147749,0.00503383482648823,-0.00299782292878914,0,-0.001799615516479
"2817",-0.0064626384237928,-0.00864787725538596,-0.00164805953911884,-0.00902356046798292,0.00505968116486466,0.00166439981016442,0.00158157408948512,-0.00375835384480216,0.00191172533127504,-0.00300482847068939
"2818",-0.00513153767813079,0.00255312095712412,0.00429188281416781,0.00161878525985704,0.0088093297779499,0.00195450786130813,0.000789871085330462,0.00653913328313815,-0.000636047071363111,0
"2819",-0.00108980246049628,0,0.00197243948870862,-0.00363624001213081,0,-0.000390167796182284,-0.000263044010749613,-0.000749421812443196,-0.00636431996096221,-0.000602764527766642
"2820",0.00108453765295602,0.00190999316278884,-0.00442923089955494,-0.00223041288364301,-0.00357623238314209,-0.00117081643468442,0.00591881837928843,-0.00248821650028264,-0.00240195352438821,0.00361883050760348
"2821",-0.0135303984910106,-0.00635444545669483,-0.0169714792549686,-0.0107700601823928,-0.00317156369166616,-0.000976872041693388,-0.00928359045057514,0.00428301152395894,0.00216697435259983,-0.0066105484132043
"2822",0.00170057479891672,-0.00127920640438173,0.00569901705385201,0.0110928675323105,-0.00401883882693832,-0.00195551037336161,-0.000791714526473752,-0.000501701837463342,-0.00448470398451106,0.00665453856253961
"2823",-0.00191921589496868,0,0.00133333407955449,0.00589171737739469,0.00109266680101627,0.000685721177630327,-0.00766103725206058,0.00175699999820145,0.0174563996051227,0.0180288471202825
"2824",-0.0249971789735494,-0.0217715806015193,-0.0091545619001514,-0.0333264468922997,0.0099095486782137,0.00411189943729395,-0.0057976907630376,-0.0122778111565018,-0.00395319408713168,-0.00767416064361603
"2825",-0.0213145688271519,-0.00654595177993356,-0.0209978389212614,-0.020267553730456,-0.000748684302117497,0.00136543438924175,-0.0159287898847859,-0.00659525167862529,0.0129385454928113,0.00892313813065582
"2826",0.0273591090406238,0.0197672985243909,0.0142417010888134,0.0324162818626172,-0.00382779859044058,-0.00272668369214291,0.012619977960638,0.011491256102617,0.0052503565139852,0.00058967534721921
"2827",-0.0170117482976895,-0.0105535320062737,0.00236844918629786,-0.0181781013925114,0.0106924899891414,0.0056627075362754,0.00270948660176229,-0.00580659295975516,-0.00615841133581552,-0.00412480965262829
"2828",-0.00295491754683208,0.00653030110832731,0.0113079615985574,-0.00504944327561785,0.00264492378389813,-0.000193887094720901,0.0193190790186464,0.00761814909446001,-0.013804965311867,-0.00414207687878376
"2829",0.0127777869295151,0.00843415779997914,0.0126836738873746,0.0209347155602471,0.00486335904281976,0.0020389851923921,0.000265165929723032,0.00856829961814642,0.000477197157149556,0.00891265673453767
"2830",-0.0215845962271126,-0.0139394327630525,-0.0201055170383647,-0.0180199716936035,0.0019731537386507,0.00101932105151081,-0.0137806677104444,-0.00849550756393036,0.0116861514294764,-0.0135452839627221
"2831",0.0128168634396764,0.00587199723548415,0.0126135557365379,0.00991363967879022,-0.00771254901366125,-0.00320020325908688,0.00658353876525219,0.00579614173714349,-0.0075436035275247,0.00537306070353027
"2832",0.0106993056109177,0.00410807521813195,0.000996530200287005,0.000417790940555385,-0.00206691847134655,-0.000583804047993075,0.0112118988084922,0.00927101828038945,0.00118760092190962,-0.00415671294288755
"2833",0.00789205084978217,0.00968996585998383,0.00497760352639665,0.00250500729323155,-0.00745760256051797,-0.00253079055176586,0.000924218554480882,-0.00099302847527305,-0.0051403243607826,0.00477048083169485
"2834",-0.0222860797189942,-0.00447854192988906,-0.0156843667246186,-0.0195749011262266,0.0109360695851843,0.00439160372438829,-0.00896757143042015,-0.0042245880270646,0.0046899521934034,-0.00712168600849572
"2835",0.00492844289350947,0.00921168873700196,0.00888968351687525,0.0010619075946352,0.00165167931164123,0.000194566592829126,-0.00173004569517299,0.0069876874082706,0.00340217583196578,0.0125522520913601
"2836",0.0159001849534364,0.0123115747977176,0.00548619125584149,0.0195203589793478,-0.00181388980453334,-0.00174869608509143,-0.0038652809775972,0.00669120463516437,0.00236558113862162,0.0171191926377148
"2837",-0.00524200527864505,-0.0067100752164525,-0.00247999544716193,0.00041624612703095,0.00355132597154539,0.000973150784383758,0.00227464097976005,-0.00147682941372496,0.00778790101192817,0.00754505613080703
"2838",0.00822692364401156,0.00654442278193357,-0.00165767266216144,-0.00041607293828172,-0.00732438620414944,-0.00359725338330574,-0.00947907224395439,-0.000246796703604613,-0.0116306142250363,-0.00403226212851959
"2839",-0.00293316402741506,0.00167765400720032,0,-0.0099895067907001,0.00232129441201523,0.000878151322297516,0.00350440779044336,-0.000739703868756214,0.00655499905492807,0.000578361080894707
"2840",0.00822174889110849,0.000628231461457851,0.00282252405627603,0.00126133853091259,0.000330880579193948,-0.000487357523468734,0.00483533907302292,-0.000493529945614246,0.00141231858954072,-0.0034682796207488
"2841",0.0106983823804703,0.00732364411588526,0.00380794051622257,0.00209944800460349,0.00272860978559297,0.00058512033903213,0.012966190974693,0.00691361400480672,0.000940241344673742,0.000580157907066337
"2842",0.000740573192133054,0.00332372089318644,0.00676232414705935,0.00858992927861801,-0.00799870174536466,-0.00389883877552544,-0.00171544708989957,0.00294264554497636,0.0007827632093933,0.0185506490623992
"2843",-0.005547700973627,-0.00434782413141011,-0.00376806615124725,-0.00581621815113909,-0.00814617311602184,-0.00274011939920416,-0.0142764637896036,-0.00537893545418178,-0.00195541653430453,-0.00398412652387103
"2844",-0.00847917183369173,-0.00270334630978419,-0.00197336088774702,-0.0125366877910921,-0.00720776337563211,-0.00333632839056919,-0.00858252237356727,-0.00147522824371837,-0.00760188883388535,-0.00171426242459438
"2845",-0.000150189589760208,-0.00125092883158706,-0.0013181751604695,-0.00804049357187142,0.000253296610904119,-0.000984790405253566,0.000676478116409251,-0.00664673000454929,-0.00797594585744166,-0.000572402055533772
"2846",-0.0134673471784226,-0.00501050401921987,-0.00362974904560409,-0.00469300176595522,-0.00455720900700762,-0.00118223800924411,0.00243320621023591,-0.0014869440669274,0.0048559145473035,-0.00515456898568611
"2847",0.00247175560500268,-0.00356705249852651,0.00314620951346956,-0.00771533191654272,-0.00669779101935153,-0.00217096978187159,-0.00215752166475558,-0.00297863741849524,-0.00649607051027323,0.00172709207715172
"2848",0.0101655598307819,0.00568545150842081,0.00610765607116259,0.0144709371328589,0.00699898864922632,0.00286756040667102,0.012162019835702,0.00896181910658189,-0.00350851595539381,0.00517234311863457
"2849",0.000938905949860791,0.00125644017985849,-0.00278913006633974,0.00617403910414338,0.00771310888875032,0.00167622932474565,0.0129507273354774,0.00542827345013741,0.00424100980842601,-0.000571629824671294
"2850",-0.00769058492884778,-0.00460064380211211,-0.00230342507559833,-0.00719417580362713,0.00176635110903223,0.00108296218984671,-0.00303165775989456,0.00147255019543868,-0.00725102788844623,0.00457659625192264
"2851",0.00177688445189061,-0.00546216725115778,-0.000824512786247178,-0.0049021024401138,-0.00360153393421425,-0.0015661924194762,0.00700665966301983,-0.00196040777034256,-0.0070631433361632,-0.00569480027258995
"2852",-0.00671754082256515,0.000422483162050957,-0.00594159518086912,-0.00792443430366074,-0.00109767085037393,0.000197364759152885,-0.00341309943423063,-0.00785665916398792,-0.000484981007881191,0
"2853",-0.00220365466108052,0.00358939538726144,0.000996147040885687,-0.00215882357228936,0.00448086979461237,0.00256466635290065,0.00039515907368326,0.00470168945845573,0.0050950019394258,0.00630014665445522
"2854",0.0129464266588737,0.00189358599307177,0.0072980290782152,0.00454350189696706,0.00151492517875185,0.00009852407142108,0.0105347386466792,-0.00123155292522592,0.00209206631873249,0.00682990607890632
"2855",0.00338331194493025,0.000840020897535654,0.00115272134924749,-0.00581532901526871,-0.00159675678256632,-0.000492189908280927,0.00547294569491719,-0.000739703868756214,0.000240878430697755,-0.000565341543789177
"2856",0,-0.00125889401430612,0.0031249413718597,0.00563248043735287,-0.0009259615985584,-0.00167358608563151,-0.00492501485908148,0.000740251435606964,0.000160520189451674,0.00282807382389816
"2857",0.00966568150258174,0.00693281568966708,-0.00852597601557492,0.00193873059813554,-0.00598198252614013,-0.0022676017272163,0.00612157741971542,-0.00271256615687376,-0.00208679676015089,0.00902412904987493
"2858",0.00935061025103212,0.00479866995352873,0.00578802364278563,0.0208558452790368,0.0080523915984354,0.00207531700904062,0.00919103620755291,0.00642936562616536,0.0068366282178618,0.00503079018948172
"2859",0.00305121866902525,0.00145341248128594,0.00756327147486946,-0.00168477017673008,0.00252223566247811,0.0000989855302335751,-0.00410481334836998,0.00147424365141879,-0.00143792938169041,-0.00611782543922279
"2860",0.000476611527864046,0.000414709517310818,0.00554834054092734,0.00126568188625709,-0.00528383663201437,-0.00216978974055426,-0.00734163946990896,0.00318932918786641,-0.00408001599999996,0.0072746624522757
"2861",-0.00688711776049145,-0.00518138237642918,-0.0102240017561085,-0.0206489608442119,-0.0113827543641416,-0.00553404045035621,-0.0147916491974689,-0.0124724996585887,-0.0161458352662196,0.00111115316920229
"2862",0.00420535001733935,-0.000833370709460213,0.00295125372881233,0.015060390314424,-0.0038378475222699,-0.00208710560058123,-0.00289735240202593,-0.00470506601162779,-0.0015512899685346,0.00554942804543024
"2863",-0.000844939538373723,0.00291906042251466,-0.000163401742595104,-0.0152608618397742,-0.00505153353179011,-0.000597097401628388,-0.00515130067213232,-0.00497661086127921,0.000572409840768451,0.00110373765033045
"2864",-0.00249997235734845,-0.00374220250275958,-0.00245255912390818,-0.00839424696747271,0.00860492379771838,0.00388587718539424,0.00225715651811664,-0.00300074809421613,0.000408654785807094,0.000551146903571942
"2865",0.0075184729282316,0.00605173579821039,0.00114737935411346,0.00607764251805576,0.00051216938931109,0.000694848936454884,0.0107297665074007,0.00652116476626596,0.000571840517217925,0.00771362090786609
"2866",-0.00278012838290553,0.00041494919300078,-0.00229218030794465,0.00345187318788587,-0.00153502692578666,-0.000396960708892169,0.00131048807017153,-0.00249207039241228,-0.000571513702526616,0.00109347875985599
"2867",0.00275120247632032,-0.0143064648831079,-0.00393821644529058,-0.000429844776896671,0.0072596559773086,0.0045644718730391,0.00850804451868825,0.00174886611267899,0.00106198019567105,0.00546159048228656
"2868",-0.00204836056892743,-0.00294484926814365,-0.00609544300093046,-0.00537745022196245,0.00796977324316694,0.00256811577393967,-0.00246602293245801,0.0017455199979941,0.00856858977828789,-0.00651827470529265
"2869",-0.00238289908052858,-0.00886084729884407,-0.00331522356708125,0.00410909005707372,0.00622494562357168,0.00394103913798682,0.0033827700908684,-0.000995660208102045,-0.00307465824337438,-0.0147621883463144
"2870",-0.0115010193121187,-0.0266070421955892,-0.0066523271469795,-0.0232610168996954,0.0219024585492607,0.0107947440365319,0.00298219433600222,-0.00971831350350905,-0.00016230013929297,-0.0094340048311472
"2871",0.0133447029749845,0.0177127259392971,0.00703177000371014,0.007938294417275,-0.00670803376347218,-0.00427173589919982,0.0126701126138729,0.0103171095682877,0.00146116565531007,0.0128852670219088
"2872",-0.00612591047716127,-0.00429738450658079,-0.00681635728959262,-0.000437554698720199,-0.001647231689475,-0.000487549813354415,-0.00178756677693193,-0.00423426240402824,-0.00218857901786706,-0.00276550571138057
"2873",0.00981796602328044,0.00820035700483768,0.00686313889643886,0.014007598951018,-0.00528339780138409,-0.00369442766209993,0.00345311779749258,-0.0002500538904181,-0.00495532095784434,-0.00665559702864238
"2874",0.00475126960499672,0.00256835230121299,0.00598498825329674,0.0101443654229791,-0.0072319915715634,-0.00353219039657782,0.00879442577410616,0.00850625094186741,-0.000979631006280179,-0.011725247698573
"2875",0.000727650642402988,-0.001708018569061,-0.00181787372697118,-0.00769225219666925,0.00234443201792778,0.00256000605008011,-0.00126341065995805,-0.000992085578002566,0.00392248907601966,0.00169489199511852
"2876",0.00836063032447187,0.010051400237888,0.00430446449222899,0.015073293610641,-0.00810290086083443,-0.0040264361844996,0.00113851213503957,0.00645603936440908,0.000569800579077073,0.00338416449252255
"2877",-0.000108361390714129,-0.00804576122426615,0,-0.0152737446793415,0.00968499028389602,0.00423986356946515,0.000631736926739457,-0.00764853820446454,-0.000488097957827893,0.00393474064972654
"2878",0.00295631837647736,0.00128084486934155,0.00296751695120978,-0.00193861551125363,-0.00300285176887438,-0.00137456033576577,0.00290433694830261,0.00198916608174371,0.00122090996890023,-0.000560017988806005
"2879",0.00133015785086643,0.010019165056689,0.00312293863799873,0,-0.00184040002907837,-0.000983349378990028,0.000251801165685128,-0.00198521715511379,0.00178848058225367,-0.000560216466350849
"2880",0.0012923767083548,-0.00654285711600167,-0.00622644970372699,-0.00259024113116391,0.00025143641901515,-0.000590518250275451,0.00503530457285839,-0.00447522211833762,-0.00332713616829172,-0.000560415101785283
"2881",-0.00319116079705728,0.00212434825197771,0.000824428753612549,-0.00670849463031409,-0.000502675669743158,-0.00118155905063377,-0.0201652129189307,-0.00174825287656166,0.00301255495847585,0.00392579808687055
"2882",0.00251799308869161,-0.000635997241210107,-0.000988485726582833,-0.00675377919983389,0.00829981546103498,0.00315477509131323,0.00997040565671159,-0.00375289260492317,0.00154229236882375,-0.0111730327424138
"2883",-0.00127590352307605,-0.00615187055271516,-0.0052770306547576,-0.00789650401000708,0.000914603792338209,0.000786452703865015,0.00101243130512008,-0.000785564839732911,-0.0165342928319248,-0.0242939171124082
"2884",-0.00205662141692353,-0.00917826376696096,-0.00729446868946304,-0.0121600608678659,-0.000913768056608255,0.000490930742437001,-0.000884974516020653,-0.00532588341018669,-0.00189545910319633,0.00868564270287542
"2885",-0.00383286549188233,-0.00844296562229896,-0.0106024591128505,-0.011038516926394,0.00581993786767576,0.00265006844673232,-0.000126544797582673,-0.00535443000142866,-0.0025596399755623,-0.0103329868542164
"2886",0.00170598205051831,-0.000222348103584458,0.000340202162659731,0.00432790510285463,-0.00876224438185713,-0.00323045045736159,0.00974573462045303,0.00281974159281484,-0.00447020684262733,-0.00116019641551013
"2887",-0.00626897511056201,-0.00778280497273565,-0.00374088028407549,-0.0140619355195974,0.0052538582847097,0.00265170209054899,0.00513907488233301,-0.00460111609617586,-0.0017462081864924,-0.0075492592332711
"2888",0.00182340714473894,0.0136708306440614,0.00494967248248801,0.0103517749528015,-0.0000829802672994706,0.000195866053957605,0.00635970278937026,0.00950181667543837,0.00241560177220479,0.0198948260359761
"2889",-0.0136130514910533,-0.0148129630723082,-0.0135869499377981,-0.0134334505239742,0.00224011893260667,0.00137129634982802,-0.00346941073778184,-0.00661430791144613,-0.00373938021403952,-0.0114746066791805
"2890",0.00221415508884304,-0.000224539087429032,0.00585386745672523,-0.00392342842006821,0.00140711281182893,0.000488842497931241,0.00395504859695972,0.00409734190998479,-0.00525479193639833,0.00986655672432346
"2891",-0.00828415385437808,-0.0096521073601743,-0.00667571799221001,-0.0192307172023261,0.00942397126669414,0.00381232031441447,-0.00537780368707241,-0.0119865883777778,-0.00570182784333684,0.00517234311863457
"2892",0.005717473759006,0.00249321517310652,0.00120625705427191,0.00850464060812772,0.000245740113544057,-0.000973812106764949,0.0106878007923354,0.00309749861242348,-0.0030359334957677,-0.000571629824671294
"2893",0.00143952569868677,0.0108522916891958,-0.00327027634511701,0.0149917639925778,-0.00343862621848945,-0.000779778453756097,0.00248826484330134,0.00720533848771754,0.00363729484319664,0.011441608389076
"2894",0.00213813459800649,-0.00715715756591695,-0.0158865502825497,-0.00992383774545491,-0.000782300612117925,-0.000684065609339202,-0.00595683074659081,-0.00715379298776975,-0.0100295236404632,-0.020927723011414
"2895",-0.0035313489197365,0.0058571705682906,-0.00122841586264011,0.000699249878264085,0.00535631102671252,0.00254270333406148,0.00749047028528871,0.00591879927639893,0.0101311340893167,-0.00115526692314427
"2896",0.008157999764838,0.0132140202181861,-0.00158117755120102,-0.00256236368294938,0.00286877605037761,0.0000973866875761953,0.0130112468537305,0.00690711884110784,0.0033712683797511,0.00578367033561245
"2897",0.00845808270533133,0.00486269973218634,0.00651070337360826,0.0137787155219131,0.00326945125602851,0.000877801670465583,0.00415886678257404,0.00685982653826867,-0.00159598484008439,0.00460028213185626
"2898",0.00900454469154344,0.00637942798680657,0.0138112053832498,0.0179682002712149,-0.00643590528223448,-0.00253363047667299,-0.00889256695776641,0.00454181517932439,0.00243985358876109,0.00515173632649257
"2899",0.00359844487216621,0.00240429284113275,-0.00379370589124894,-0.00226303920589843,-0.0000820878882533682,-0.000781557218396456,0.00307284331683122,-0.00276307776301643,-0.00184642884017738,-0.00227787321992068
"2900",-0.00731452594293713,-0.0183165307738747,-0.0138481548306009,-0.0195053850038494,0.00385412943704244,0.00205335334036572,-0.00306342987680763,-0.0130981942351691,-0.0108467249642648,-0.0348174624831071
"2901",0.00906591086638087,0.00888486545947265,0.00105321151922144,0.0136478616071405,-0.0000815213508297274,-0.000390446049809867,0.00294991471911499,0.00535989641536494,0.00416523294938154,0.00532240485517366
"2902",0.000787504230135294,0.00286217306127057,0.00929340685318625,0.000684569130120716,0.00253234080826159,0.00165935775843673,-0.00343120209214609,0.000507484532478397,-0.00440189632782273,0.00176480282097224
"2903",-0.000894029110107386,0.000438968253788863,0.000347544309366787,-0.0054731454420025,-0.00415574101703808,-0.00165660885168595,-0.00455012955810019,-0.00050722712255924,-0.00051014369092639,-0.0211392979429703
"2904",0.00404506745696809,-0.00175526563384854,0.00885708552374198,0.00733780919417737,-0.00188197011205604,-0.000585729496751064,-0.00531183494262721,0.00025375704189079,-0.0108039469807585,0.00119974367765274
"2905",0.00210390903204294,0.00241794110338645,-0.00154925913017978,-0.00113813184863587,-0.00401719138749423,-0.000781328285443861,-0.00471925350665403,-0.000761432522448424,0.000257989338303899,0.00898741846514817
"2906",-0.00377161362019207,-0.00350887312769266,0.000172373094012412,-0.0123063376474055,0.00633822448643917,0.00273710403535121,0.0101071529335934,-0.00558788648981534,-0.00429885657809059,-0.00118763226939633
"2907",-0.00114293335928239,0.00572192067281829,0.00310286308121221,0.014305446986435,-0.0122689941551291,-0.00350943757628619,-0.00840024167587727,0.0109835278004751,0.00647612479882786,0.00713438888152895
"2908",0.00185923578325498,-0.0026257918121444,0.00498369717082081,-0.00659697407977156,-0.0123385583261743,-0.00489157344821889,-0.0024915671112441,-0.00480053252263646,-0.00480437551139967,0.00354192497063477
"2909",0.00503221966219991,0.00680103166609403,0.00410406706379352,0.014655431755308,0.00343761621287197,0.000688172624575545,-0.0048708877457786,0.00330026000714256,0.000344836206896515,0.00529404521019172
"2910",0.00852248844185177,0.00740920767367204,0.00647126278708687,0.0162489548490226,-0.00158787777029201,-0.00068769936869606,0.00815797723764344,0.00607284575531408,0.00551533087284284,0.0134581601662647
"2911",-0.00235895822717402,-0.00605656079584671,0.00253817696186354,-0.0111035795189581,-0.0019246695744306,-0.00108145375495994,0.00273851347380338,-0.00829974511461873,-0.00779913438464175,0
"2912",-0.00677654353154999,0.0019585885743354,0.00303797809173822,0.00359309255454177,0.00167694832494547,0.00157465276736701,-0.00968340215794072,0.00152188340629,0.000518312184114356,-0.00404145601756001
"2913",-0.00522353067917403,0.00260640046778682,-0.00757202068340912,-0.00156638261294406,-0.00343188476836942,-0.00127719430704909,0.00137877463805136,0.00177244940209786,-0.001554001527169,0.0057971412257396
"2914",0.0049293619864188,0.00411595188041569,-0.00762965239587299,0.00537876790198633,0.00545972143402773,0.0013774386394978,0.0171508169312911,0.0045500875373321,0.002939870247473,-0.00576372808007275
"2915",-0.00167040197624191,-0.00755108437756191,0.0064924124571768,-0.00891658157573461,-0.00814689378723132,-0.00236289562790881,0.00332319356554578,-0.00603957740415628,-0.00732820945474966,-0.0144927933996526
"2916",0.00544749672025202,-0.00913043833423566,-0.00560166277654939,-0.0132703621797172,0.00143504620495905,0.0011840504992866,-0.003312186528586,-0.00278452741053248,-0.00538476641814112,0.00588239354001052
"2917",0.00428483723550999,0.00197451109390379,-0.000170808620166718,0.00775019672331068,0.00497361922773365,0.00256272057490969,0.0118155143404444,0.00406197440236533,0.00349284850225762,0.00350872377936784
"2918",0.00366707357198237,-0.00459829946452572,-0.00751229404568843,-0.00769059311376008,0.000587135995162358,0.000491637774077347,-0.000608090867361799,-0.00455135561179631,-0.00513397154775463,0.00174822784108608
"2919",0.0033025217543412,0.00791919732121604,0.00842921911704497,0.0102575841312766,-0.00519765829215857,-0.00206353804740844,-0.00352975647015885,0.00330184825861335,0.00227406625952842,0.00756249299486456
"2920",-0.000420268196043683,-0.00174587377098412,-0.00102344203448057,-0.00135381201444873,0.00101147876580421,0.000886391432732614,-0.00598531809338021,-0.000759151345356535,0.00279263470783264,-0.0121246057469363
"2921",-0.00136605555892677,-0.00349813283464295,-0.00375692172155384,-0.00293715188581478,0.00841808710346137,0.00275451883086575,0.00122878490031764,-0.00354713776473559,-0.00147947083876176,-0.00409111864171874
"2922",-0.00670038844313781,-0.0223781184320072,-0.0143982944895316,-0.0213007020829639,0.00726266754192118,0.00431646243734884,-0.00895903479649574,-0.0142383190530269,-0.000435732969073177,0
"2923",-0.00374318792298578,-0.00269313505923674,-0.00591304219955291,-0.0164389428758146,-0.00207185815447708,-0.000292993511806228,-0.000495335208985925,-0.00464313259048665,-0.0150841657496876,-0.00528167780563416
"2924",0.00638064780660841,-0.00180018416734118,0.00402386324938653,0.00612057368480423,-0.00224247933852417,-0.000977145312029415,0.0054516551479824,-0.00259117229589978,0.000973804895306296,0.00176976566726261
"2925",-0.00746742952840429,-0.0171326273025196,-0.0121972700817402,-0.0287788526245893,0.00582673227988506,0.00244524754610342,0.0075169035386291,-0.00545586132431675,-0.0166268506235074,-0.0217903474683254
"2926",0.00809129893596827,0.00711025173830548,0.00546836807796902,0.00626377836630732,-0.0000827334757773635,-0.000292803101282435,0.00807235143361118,0.0070532728526429,-0.000809461267929579,0.00782656574689478
"2927",0.0035205216352483,0.00592110082029218,0.00333324046776839,0.0105337360629847,0.00124135702162453,0.000390599922918566,0.00897841261217458,0.00648493752049695,0.00927091825870252,0.00418166710267975
"2928",0.00214020243077573,0.00701832754220266,0.00402166148146899,0.00450136158209391,0.006695272376122,0.00312180862308731,0.00156328651022464,0.00670124983994635,0.00499424788176883,0.00178462762613107
"2929",0.00234513971506645,0.0107913682799481,-0.000174114244333334,0.0127358242921018,-0.00336654540734482,-0.00136150149202341,-0.00672335607698127,0.00179196195203257,0.00292834319055202,0.00178144840409455
"2930",-0.00059362840457311,0.00333637460718506,0.00418041275399905,0.00791795226564185,0.0039547349971738,0.00185039887924443,-0.00556041973975763,0.00178887555896212,0.00221199793519733,0.0142265489565536
"2931",-0.00132799344853718,-0.00753729557224703,-0.00416300965534089,-0.0161736406692967,0.00155888195452669,-0.0000970174161267767,-0.00218816057205573,-0.00612245007041168,-0.00944645562231283,-0.00175333656073662
"2932",0.00601829080943195,0.00826454510741659,0.00348372566345123,0.0185533664384234,0.00196674524050633,0.000291526681871046,0.00511662836935622,0.00487692830272146,0.0174688685597737,0.00761113664734459
"2933",0.00789531208522187,0.0132921410167444,0.0151014684817035,0.0142955509081295,-0.00572416107368712,-0.00223558953100145,-0.00181804528120555,0.00791823002423153,0.00376657309857831,0.00348629761126173
"2934",0.000483316858928218,-0.00174911283073864,-0.0030779968789475,-0.00363719919011829,-0.00600391482106699,-0.00224013120568189,0.0106847692942638,0.0012671834674105,-0.00794132150942739,-0.00405309730294123
"2935",0.00538070126241563,0.00459912036133292,0.00360211928328202,0.00616005530910813,0.00132376884771679,-0.000292903272347544,-0.000961023100099268,0.00556808538852449,0.00457421710063333,0.0110464194354272
"2936",-0.0040482146574673,-0.00981025560768101,-0.00700735039081612,-0.0260770892909589,0.00214869625118297,0.00185514257989183,-0.00348731146884285,-0.0113264440264668,-0.00490366037400147,-0.00172510579944607
"2937",0.0000343960179549629,-0.0112286383421585,0.00206545467110941,0.00512226681259054,-0.00230882591403925,0.000195174500603912,0.00374089270941402,-0.0015274580468374,-0.00114393700408255,0.0011520579548232
"2938",-0.00172225244920865,-0.00823861600478459,-0.0123669158810873,-0.019457944662461,-0.00578147956726272,-0.00228512711639051,-0.0105794367204913,-0.0114736089779459,-0.00510969949590867,-0.00575372044135014
"2939",-0.00269154007348271,-0.00583744513885431,-0.0106087088045981,-0.0144105226088038,-0.00266616744542025,-0.0000976286537959226,0.00461707931365019,-0.00438510738820364,0.00345346674931357,-0.00405098955429095
"2940",-0.00300996066685688,-0.00496831660183794,0.00228513968777544,0.000958584293588638,0.00367567647860101,0.0020552522287709,0.00387044249218937,-0.00103613396190749,0.00194141369572898,-0.00581049601876982
"2941",-0.00194346967428372,-0.00817065856881294,-0.00613817260976834,-0.00502852332555714,-0.00848943751950526,-0.00449324900685155,-0.012168680648961,-0.00674280712148367,-0.00273029766839628,0.00233778208098223
"2942",0.00173848468224791,0.00892447768876936,0.00229393726382932,-0.00986772040758821,0.00369343089051322,0.00058862485456368,0.00634231289100962,0.00104446257042579,-0.000706535351765347,0.00349849440394534
"2943",0.00329740518206423,0.000453504257516002,0.0021126540438714,0.00218762195904709,-0.00761062729401385,-0.003628420606413,-0.00206047574845947,0.00365159229875123,0.000618638963877371,0.00987802264203652
"2944",0.000242379412822347,0.00385403748664848,0.00193253814414751,0.00509334333193268,0.0023596956351366,0.00118091347028337,0.000850061856658701,0.00545727852820677,0.00839071711366635,0.00690439346752192
"2945",0.00591432872323838,0.00722675565157527,0.00771529735310383,0.0135136765565944,0.00151353097965168,-0.0000983778089791443,0.00594602111613063,0.00361852911468374,-0.00359110105266014,-0.0108571717928199
"2946",0.000171893893074593,-0.00224213976597953,0.0113102785186934,-0.000952370625918797,-0.00478529248042669,-0.00186812385909074,-0.00808210695072609,-0.00309043932730046,-0.00650496648198018,-0.00635450319835917
"2947",-0.00529428586439584,0.00269669500590108,0.000516087396412956,-0.0090563860906191,0,0.000197143264285105,0.00352664726029062,0.00258313929893594,0.00522035051903247,-0.00116289437072703
"2948",0.0054263320484027,0.00515450490106639,0.0239036964260244,0.00961995765157875,-0.0104599694063963,-0.00413615795245492,-0.00351425372701231,0.00669973388760292,-0.00149633833732643,0.00931320734642194
"2949",0.00106552604287802,0.00222973656603953,0.00352703019660638,0.0138161705860607,-0.00596684301507355,-0.00168124438644535,-0.0132555607514251,-0.00358357233548057,0.00387865825319711,0.0063436269774495
"2950",0.00810398941424095,0.0180199008013298,0.00267781968258807,0.0110432206468689,0.00463077983203797,0.0000989631922199141,0.00998277687056248,0.00796306787491363,0.00342465762446409,0
"2951",-0.00091378706486922,0.000437139370168316,0.00216993087935058,0.00464804295070742,-0.000426615032298128,0.000396081680468674,-0.000487871212014435,-0.00790015837753066,-0.00682592999455489,0.00229223237918608
"2952",-0.00332196388582962,-0.00480552772024068,-0.00449694658220268,-0.0113347150840254,-0.00256203615707873,-0.00108892220500068,-0.0175804001125583,-0.00363341751416846,-0.000176200549408811,0.0148657296621684
"2953",-0.00092774133535789,0.00570673237435582,0.00752882550862144,0.00397741476360736,-0.0010272834458247,-0.000991252288833899,-0.00161555842126015,0.000520875315407565,0.00158633117488027,0.00225360625707682
"2954",-0.00299215033893452,-0.00152767140312604,0.00481568045524194,0.00209735978716519,0.00702766734772786,0.00327430599031064,-0.00915046055595903,0.00364488888474312,-0.00527935758417319,-0.00449707787132436
"2955",0.00279394939351363,-0.00284162049792236,-0.00264418643555353,0.00488371204873217,0.000680775630213182,0,0.00266390657074211,-0.00181584090100562,-0.00884564328582993,0.0045173929391471
"2956",0.000103465184353224,-0.0120561175442319,-0.00198838026586334,-0.00671150370612372,-0.00263668126992467,0.000494581138530625,0.0123986076111338,-0.00597714951804718,0.00633644784462883,0.0101179045278676
"2957",0.0034742361713811,-0.00044371397547105,0.00680723985039067,0.000233131365295236,-0.00734087832461716,-0.00253570428068184,-0.00824783426899367,-0.00261436105271873,-0.0016850123858636,0.018920451388869
"2958",-0.000582987242476962,-0.00532733189612045,-0.00230876314268258,-0.0125785682977757,0.00611238052700847,0.0025818965058817,-0.00138586901379223,-0.00996076362965514,0.0115483965532557,0.0032769655314917
"2959",0.00054879740873659,0.00379364151684269,-0.0087603112728758,-0.00825665694092736,-0.0173710507374152,-0.00742799778731817,-0.00694018943286789,-0.00529514115536756,-0.00395191875071776,0.00925425988695894
"2960",-0.00781576585140542,-0.0131168861939245,-0.0135067950969243,-0.0249762916628088,-0.00705403713121977,-0.00259451956902057,-0.0100382752954604,-0.0188980492309569,0.000529051323030272,-0.0107876155675189
"2961",-0.00559694293234547,-0.00698354400546652,0.000169010842832273,-0.00365939653468317,-0.00859492059233735,-0.00240105750210851,-0.00128337259419975,-0.00189912698355899,0.00281988008054612,-0.00218110757682066
"2962",0,-0.00930131878631035,0.00439422570538706,0.00146927511974537,-0.0033614839926247,0.000401552657775195,0.0132372289238669,0.0046209770739527,-0.0110720735218258,-0.00273220340393854
"2963",-0.00145933248552832,-0.00114501724744964,-0.00572108501972313,-0.00366755222786652,0.0101188921777453,0.00190421433455157,0.00215630272552891,0.00865769857118615,0.000533117109177805,0.00712324725195068
"2964",-0.0316630291597867,-0.0194863171190136,-0.0245388633052572,-0.0296932379686408,-0.0027241643770719,0.00050030761736175,-0.015061357403946,-0.0179719206779069,0.00248666967116651,-0.0195864096426023
"2965",-0.0220266541106497,-0.0126257191324982,-0.0180429953621853,-0.0101163899230214,0.0121598630488828,0.00410015098858896,-0.027242342941638,-0.00409721295427967,0.0256910176920009,-0.0149833186461571
"2966",0.0138883944266042,0.00189446762167078,0.00229677446322363,0.0293817780105878,-0.00348225820997894,-0.00119510682548274,-0.00198137930618492,-0.00191989894683298,-0.00475035416091174,0.00788721601174891
"2967",-0.00561700519768482,0.00165443064529902,-0.00299654944348804,-0.0106726992780348,-0.000437093497130392,0.000598118204524045,0.00542661080003404,-0.0010990055035438,0.00668226138985695,0.00223597067338011
"2968",0.0218657509658873,0.0160452025003821,0.0185643558432182,0.025087911245947,0.00227253059737564,-0.0000994473332988077,0.0217221361123712,0.01980734992445,-0.0017241120689655,0.00446184972113572
"2969",0.000178392877584699,-0.00952147518501423,-0.000694268449732194,-0.0122370468870082,-0.00592953832918897,-0.00289008860617801,-0.00489636911984825,0.00161848590733493,-0.0000863730547572272,-0.0088840601011867
"2970",-0.0144411778296949,-0.0164128157175335,-0.0180650580849466,-0.0262635704626462,-0.000350828328708142,0.00179903246867541,-0.00116537829414209,-0.00430921592047417,0.00112269625077555,-0.0112045023045214
"2971",-0.000542353273061624,0.00786647893951287,0.00212274458617978,0.00941475847591078,-0.0021938068832511,-0.00119725300042672,0.00764866496892869,0.00405731559710931,0.000776432035480168,0.00566582033804575
"2972",-0.00448881433969783,-0.00591292831448109,-0.006178263412287,0.0108394226006892,-0.00131915239221736,0.000199444088647915,-0.0131224854175576,-0.00484919747850288,-0.00258600978215662,0.00112674514453537
"2973",-0.00509076075286563,-0.00713769354177674,-0.0115451944998513,-0.0109725037383912,0.00316996524966973,0.00259676943008014,0.00638765825286036,-0.00378981004948209,0.00587676091847511,-0.0219470914597191
"2974",-0.0302986453198093,-0.028277001266317,-0.0319856688491623,-0.0322743847446737,0.00754930570468981,0.00537905800839122,0.0072538279636496,-0.0138587867377079,0.00231982990222379,-0.00690445268593698
"2975",0.0179406831378834,0.0128236382801217,0.0148505396962857,0.0192807374231192,-0.00418180490328535,-0.00237774489327236,0.0123457655968211,0.00909341501222682,-0.0022287158502069,0.00405556430793319
"2976",-0.0175874435884369,-0.00413920969194115,-0.0128041033838174,-0.0115029657898348,0.00603660211205526,0.00446910779573506,-0.023500990310543,0.00191163642766612,0.00317865114813309,0.0075013995081854
"2977",-0.00554018645677168,0.000244424713295333,-0.00926434169429746,-0.0173261059878479,-0.00226084696535467,-0.0000988965190500402,0.0115778754116609,-0.0032708742507922,-0.003939359525718,-0.0103091969184586
"2978",0.0148182188719781,0.00855539506148184,0.0157096763030147,0.0194738809173298,-0.00496833466707569,-0.00217530169965774,0.0150464387786904,0.00464896563727879,-0.00438479072108655,-0.0052083811063095
"2979",0.0106811010815482,0.00799813410915506,0.009758770252144,0.0108413482972176,-0.00508060042479885,-0.0024774920762175,-0.0103888774357244,-0.00816558587094796,-0.00561313456960799,-0.0133799887343048
"2980",0.0106419194879068,0.0158691899499488,-0.00237054260309932,0.0357508160388309,0.000926868430329852,0.000855992023635066,0.00371276346120109,0.0148187763431475,0.0128527570498871,-0.00707537594761776
"2981",-0.00592315614836414,0,0.00566625423388833,0.00641009568806217,-0.01243293208313,-0.00557041405133718,-0.00854595073654207,-0.00459704770842029,0.000171525340946443,-0.00237526453879289
"2982",0.0055170199478658,0.000709894312775683,-0.0036350544341196,0.00269481336195332,0.00392867021048415,0.00059992738114123,0.0146660984493461,-0.00135831710394774,-0.00240033429232178,-0.000595229963322619
"2983",0.00632782408344079,0.00165568018207951,0.0113097310259052,-0.00171009553395529,-0.00062271222773469,-0.00109934560027902,0.00431097785114343,0.00788895490527697,-0.00283579953160262,-0.00416921391002356
"2984",0.0214088704754858,0.0129870904586253,0.0104618646677477,0.0188447814972832,0.00133491097847593,0,0.0126243363999243,0.0156546927075201,-0.0000861944149759264,-0.00239218884047798
"2985",-0.00181500179084881,-0.011421965187482,-0.00642628327143213,-0.025942958349894,-0.0000888797526600316,-0.00140126062931034,0.000374098338149498,-0.0087697203976933,-0.00215461520429727,-0.00599530645430091
"2986",-0.0097680201251239,-0.00377260377338462,-0.0100611231213116,-0.0184957297892748,0.00746626603190581,0.00390870949346289,0.00137117650782437,-0.00482576550211766,-0.0112281569461752,-0.0108564294470516
"2987",-0.0186853796404133,-0.0201182782007877,-0.0136116904106344,-0.0140702027728276,0.00652833187078472,0.00299498270360465,-0.0011203258316671,-0.00592668311857114,-0.00716281427770404,-0.00243899102184708
"2988",-0.00187085016844035,0.00748770496784057,-0.00367978910579181,0.0114678952442575,-0.00061377956668629,0.000796255893785514,0.000872343323208735,0.00785914875831506,0.000351865199652801,-0.0275061756106754
"2989",-0.006836685704109,0.00119874660943831,0.00350875135019635,0.00604687845268548,0.000614156523411014,0.00208844816335829,-0.00174297964350845,0.00349538385361603,0.00826738808093386,0.00879950644204519
"2990",0.0104365830913273,0,0.00588891443304318,0.0222888656189077,-0.000438127802642962,0.000694825435847868,-0.00623517513709004,-0.00535898920978606,0.00113396721156644,-0.00186913334812067
"2991",0.00260051910881964,0.000239518187928001,0.000731661888079715,0.00196003684310675,0.005787308064515,0.00307443786594108,0.0120466567454001,0.00377168080218038,0.00740616905304958,0.0062422403245177
"2992",-0.0169145791562346,-0.00766094236770121,-0.00438752317372226,-0.0134475530791679,0.00278981344011431,0.00148289869123786,0,-0.00214715223356643,0.000432407876689078,0
"2993",-0.0185060975345984,-0.0176115466757807,-0.0183620309598644,-0.0215612980160856,0.000347773516385264,-0.000197321986527554,-0.0106633849356863,-0.0134481825295959,0,-0.0303970519984572
"2994",0.00340753088259538,0.0135068771817486,0.0153384948608142,0.0184903037241231,-0.000347652612013971,-0.000197432586117929,0.00137870859545441,0.0111779279267255,0.00164262992379394,0.00831735623043794
"2995",-0.00667878971264857,-0.00799609278468671,-0.00368461127184183,-0.0116884371725613,0.00104352923141193,0.000592496628997408,-0.00337922464811635,0.00242645083001669,-0.000776834103427881,-0.0291878088056222
"2996",0.0161444877911301,0.0158768794930704,0.0134985892990058,0.0123299516319388,-0.00225837985336785,-0.000789735774091249,0.00351618726434966,0.00968258854723381,-0.00112289888026862,0.0045751006142738
"2997",0.0033644161785038,-0.00456834902907322,-0.000912235934427907,0.00696001123645584,0.00113178217548082,0.000988024181436398,0.00312867205272194,-0.000799111344238712,-0.00596681084371165,-0.00390365519694513
"2998",0.0230252456048836,0.0132848189767496,0.0131482411501289,0.0239447823299515,-0.0048693335591895,-0.0000987345637727399,0.00885721522813032,0.0130633070698596,0.00374075694843223,-0.00326592898342237
"2999",-0.00218506996109036,-0.00452922164881775,-0.00342463754381817,-0.00867891561743406,0.00393187834704234,0.00256615505769076,0.00136019035022117,-0.0115789864939716,0.00312013355313234,0.00655312555937493
"3000",0.00609534065601314,-0.00574703849473879,0.000904316374224612,-0.000972674727714673,0.00374241085987514,0.00196869858143867,0.00987884792801874,-0.0106497361690016,-0.00172798516896466,-0.00455729637804392
"3001",0.0132412367288259,0.0108381656393342,0.0135525086914956,0.0202043179263898,0.00710026731013191,0.00218599339472969,0.00464679308357097,0.00188363987293294,0.00752988568868029,0.0228908020595362
"3002",-0.032402310650007,-0.0228734321746841,-0.0369048430383533,-0.021235849728057,0.0167416361071027,0.00461729925667909,-0.015457819438196,-0.010475289518048,0.00609912357704245,0.000639377437478439
"3003",-0.00151695287134879,-0.0141429818338963,-0.00148096887147153,-0.00926389340754274,0.00314033820817361,0.00254236884339143,0.0250958657784317,0.0114007283219246,0.00017073086994368,-0.00830666140199077
"3004",-0.0232361098518953,-0.00964629515951909,-0.00741553739108447,-0.0187006916097683,0.00186165298508945,0.00292614876199848,-0.0141100151412102,-0.00161038736490116,0.00810992836016666,0.0115979115668692
"3005",0.00189707896627644,-0.00774213983602179,-0.00765796228353266,-0.010531733842116,0.00413814253895772,0.000583461911908056,-0.00562690428753221,-0.0083335230215712,-0.00347189443549467,-0.0159236109303792
"3006",0.000227130022296906,0.00352362632515368,-0.000752810210529087,0.00760267554393335,-0.00016835711035279,-0.00252672655290442,0.000738256237766688,0.00135546536608455,-0.00118965839564922,0.00582522978331501
"3007",0.00503538321253627,0.0175571218398687,0.0120549792476998,0.0163480937218123,-0.00445822092345671,-0.00272879644835389,-0.0164719928406142,0.00730909982304206,0.00212693549321985,-0.00321752554992527
"3008",-0.000338944551161791,-0.00172549205526418,-0.00297792445084577,-0.000247401743181497,-0.00236601785218116,0.000586350046671624,0.00599907691087997,-0.00322470083750004,-0.00220733506912862,0.0129115793058858
"3009",-0.0184647984097039,-0.0143209758504466,-0.0113869849133919,-0.0141089362560833,0.00347277042660687,0.00156248516193225,-0.00198763025257431,-0.00350502527664254,-0.00399898752658046,-0.0152963551974954
"3010",-0.0196183179190484,-0.00926844267678484,-0.00793041170494901,-0.00928956035297224,0.00582356722094324,0.00292524939725847,-0.0369156901220846,-0.00730520591225381,0.00691957127831144,-0.01165045956663
"3011",-0.00109653752344296,0.000407466814616564,0.0027812194198753,0.00679092397450898,0.00598882387574773,0.00246468035400049,0.00897151581944988,0.00109020768362167,0.00237548988609082,-0.0209561733922374
"3012",-0.0149757176260689,-0.00687367808981643,-0.0147283493004392,-0.0166070454245462,0.0132107438979046,0.00349854043132902,-0.0109535169352218,-0.00490074874231783,-0.00609396519519312,0.00401346090748089
"3013",-0.0162779530052772,-0.00410155002733237,-0.0052417117512894,0.00779417915395775,-0.00363101221313122,-0.00125916142764226,-0.0145929991377908,0.00136797965606217,0.0154134207613046,-0.0093271930529496
"3014",-0.0204895671992901,-0.0123552718203471,-0.0308353416759635,-0.00696057448498988,-0.000165726076835515,0.000873012515615113,-0.0124287471128718,-0.0191256462506961,-0.00436092761423901,-0.00874238444107645
"3015",-0.0264230088264695,-0.0125096419736017,-0.0108738833895117,-0.00934589969424127,0.00497036927341554,0.00251868835736491,-0.0360156106093414,-0.00725830325740995,0.0109501009859325,-0.0110645613123692
"3016",0.0505249907638932,0.0250724893552119,0.0189331879385217,0.0199162076833277,-0.0107154634762509,-0.00473526646284184,0.0327778036156825,0.0187104439739849,-0.00299944183468026,0.0222376880571071
"3017",0.00767733058360931,-0.00411939391576455,0.013386713485267,-0.00128459731383579,0.000166460614608566,0.00252477489937286,0.00161368145461749,-0.00367344112695389,0.00760484681247364,-0.00951735773123952
"3018",-0.00128999284734821,0.00853152183069406,0.00118281834727685,0.00951885530401997,0.00841400824113747,0.00542343865768125,0.00308822650789065,0.00226894572547165,0.00406401260678435,-0.00823610138714159
"3019",0.00875885574148416,0.00281962148382031,-0.00177227384930445,-0.00458711439609583,0.00379994724488375,0.00375709335346719,0.00307849106384728,0,0.00156948623111663,0.00276814258750346
"3020",0.00104026095597276,-0.00536801862746317,0.00690472741629278,0.00256017326894109,0.00526727776148839,0.00211108700080809,-0.0216173238638049,0,0.000659810309278308,0.00276057124542151
"3021",-0.0238628403463345,-0.00719597733110466,-0.00568183474559802,-0.0181308682721302,0.011379198598936,0.0079488102005334,0.00641011067965525,0,0.00906616650348369,0.00825877456338286
"3022",0.0334958416311826,0.0300283881935774,0.0338916189680742,0.0322496993501982,-0.0115748569827321,-0.00807598016857847,0.0107061883101598,0.0209394651155193,-0.00808623703340683,0.0136518996195234
"3023",0.007884650261337,0.00150786756751531,0.00247752185742289,0.00226765866061429,-0.00294833295373664,-0.00277795513829249,0.0100565393839813,0.002771684274254,0.00345848973223828,0.00740742970686781
"3024",0.00939525742480041,0.00727732259179259,0.00475293652472142,0.00377076610839233,-0.00262834882310892,-0.00249731638169615,0.0181861984974756,0.00801551230077258,-0.00270804199320496,0.0100266691442319
"3025",0.00467351978092601,0.0122073725401903,0.00548716592059284,0.0177810536769176,-0.00156478422687922,0.000577850592822005,-0.00130369294522525,0.00740321191470494,0.00641816017788321,0.0198544006138881
"3026",0.00352751342297219,0.00147669322388833,0.00602185322959459,0.00713592795280493,-0.00643340649017587,-0.000481027275638479,0.0138382837872988,0.00653239187907984,-0.0058866978315214,-0.00259576096476599
"3027",0.00038634581348318,-0.00466950295466462,-0.0115973439267836,-0.00488651129763962,0.00390165767312567,0.00298465525328839,0.00347673009585359,0.00216335247084953,0.00172717334409644,-0.00325304643822777
"3028",-0.00610081946632579,-0.00419739889597759,-0.00359569218570532,-0.00834756840673112,-0.00372108834094953,-0.000576144794930844,-0.00320815117902262,-0.000270020909575508,0.00238089485104531,-0.00848568371229008
"3029",0.0114607621218774,0.00223145130274305,0.0121555561220799,0.00693227380274131,-0.00365223783475677,-0.000960196616154985,0.00991247365206238,0,-0.00172003445720481,0.00790000123072776
"3030",0.00241972641519861,0.000247442040853807,0.00487905024293855,0.0122941465384012,0.000999765623281634,-0.000577100471074954,0.00624608582167596,0.00296912270604754,0.00319986880209711,0.00522536480298497
"3031",0.00758683582852049,0.00519408512986552,-0.00205424078648098,0.00437205057862333,0.000249564267445157,-0.00182764129666679,0.00532055905030604,0.00376752086229781,-0.00130854669113967,0.00064975053065397
"3032",0.0133100443457361,0.0125493890557979,0.0132859550808924,0.00483687882741157,-0.00524152109106435,-0.0031804019994458,0.00378038750730081,0.002948981002872,-0.00892641054027998,0.0103896539161537
"3033",-0.0135105694448745,-0.0133658840692076,-0.0179131622341139,-0.0173284876704741,0.00677475176448272,0.00348037322047867,-0.00288740969138102,-0.00534620117490536,0.0035531318018458,-0.00706942989049986
"3034",0.00209240277831846,0.00689664802852485,-0.00282062818466799,0.0102864940062133,-0.000415165892432845,-0.000481722734633538,0,0.00618128128818141,-0.00139973655166081,-0.00129445445557619
"3035",0.000531402569220463,0,0.00584569091438558,0.00969703082132423,0.006565774557592,0.00318117502916127,0.00352505946020076,0.000801151041986747,-0.00156664744035828,0.00259226447945782
"3036",0.00846157782732559,0.0102739217532575,0.0108735957904251,0.0132052421422242,-0.00478913397522429,-0.00230603965880727,0.0116673183948024,0.0122765702015997,0.014617268630515,0.00517138674472584
"3037",-0.0076002856358115,-0.00460053462569421,-0.00723288362161978,-0.0104266380048906,-0.000995640715207413,0.000288936135260931,0.00905248131945835,0.0058000884892242,0.00349991857805709,-0.0135048870193266
"3038",-0.00132704448333043,0.00316237145047715,0.000934049132038206,0.0016764193165979,0.00506609124680146,0.00288841741426182,0.00798819056842737,0.0104848829323478,0.00559657713037076,0.00977835680421557
"3039",0.0158309237536634,0.0106691782039003,0.011198245690329,0.0217547021442757,-0.000743758562761432,0.00230411645283546,0.0079248850762057,0.00804146311416098,0.00572672191337187,0.00710137726681648
"3040",0.00878238431921341,-0.00143959369876701,0.00184562933137644,0.00842292121598209,0.00860004998328168,0.00459764929752438,0.0105238918189394,-0.00205872129710782,0.000481177312035008,-0.00512816137458549
"3041",0.000481601871410442,0.00120136139099269,-0.00405292340605612,-0.00788864581837989,-0.00603968496400964,-0.00535063787014955,-0.00682306046164505,-0.00128923940174619,-0.00200400801603207,0.00902057392904099
"3042",0.00703535362097729,0.00287992903660617,0.00221969038213921,0.00163711610463801,-0.0044642261216099,-0.00220925722558107,0.00674930565095466,0.00206563146751204,-0.00433735742971886,0.000638547936024469
"3043",0.00419200053884361,0.00909288033612432,0.00406053709978149,0.0137753413215211,0.00456723537454518,0.00173281516196244,0.00610575925330825,0.00154620368597524,0.00258147791692065,-0.00446711284627554
"3044",-0.00131831329145282,-0.00450542246763286,-0.0082720766655241,-0.0135881597825848,0.000496039357047673,0.000768528444364369,-0.00690154618172245,-0.0061744286865838,-0.00675890736046758,0.00128200777892928
"3045",-0.0095326937110336,-0.0131015229905782,-0.0139017208981284,-0.0100396625750961,0.00660981688619122,0.00326548378201097,0.00766822951892943,-0.00310638001972363,0.00243029808116813,-0.00960307277514072
"3046",0.00122148091037322,-0.00362056152965529,-0.0088345902156145,-0.00566048174513201,0.00426827847051614,0.00133984813187471,0.000237914858662647,-0.00103877404483266,0.00379829487309347,0.00129284668618146
"3047",0.000554537745337091,-0.00242246139988722,0.000948082963588615,-0.00332065581122831,-0.00392300529811329,-0.00152934116097814,0.0028530986852624,-0.00285938016550047,-0.00491104584905433,-0.00581019987504727
"3048",0.0128593803973338,0.0109275734524532,0.0176204161877671,0.00832931070506926,-0.00254373047928691,-0.00134018372234235,-0.00580850372152764,-0.00052153514183706,0.00210358417643342,0.00584415558710938
"3049",0.00324677932409378,0,0.00242040046765846,-0.00708040935766341,-0.0037842628068131,-0.00249264210937949,0.00465011012411387,-0.00756381843660692,-0.00395606326533127,0.00581019987504727
"3050",-0.00221798795341488,0.000240249991621422,-0.000743009777828374,0.00190161948145717,0.00569785835938585,0.00470918967624989,0.00320440131503719,-0.00289109012230748,0.00559289116658279,0.0025673722456947
"3051",0.0108970914385698,0.0158500335639045,0.012825378107119,-0.00142343320556615,0.00156001098711456,-0.000956566788778423,0.00615162729165597,0.00711649212989895,0.00596489611421736,0.0185659623806202
"3052",0.0017306129349226,0.00401908537407469,0.00165175861519495,0.00784020391447648,0.00254131794392953,0.00172351617975486,0.000235157351440751,0.0036641086404452,0.0152243105314669,0.00251418451559937
"3053",0.00201548493278403,0.00565088848131956,0.00109922401747409,0.00565771500944212,-0.00286197401731536,-0.000191277343502438,-0.00705299948323523,-0.00260774098544003,-0.00173633784695348,0.00313475350515446
"3054",-0.00355581707206409,-0.00468273206620007,-0.00146412989547584,-0.00210968555668289,-0.00893878057770381,-0.00296369665132057,0.000828513291079025,-0.000522682813473674,-0.0113061350891966,0.00312495753357278
"3055",0.00619992593121754,0.0030581989638212,0.00219942454183175,0.0110406726155554,0.00595779945507724,0.00297250625816403,0.00532318661072817,0.003138882531734,0.00359853649903541,0.00249225404025921
"3056",0.00136127853545021,0.00211066259023052,0.00566942618248123,0.0111524039816433,-0.00296125715129625,-0.00152956601046361,-0.00729506112415612,0.00104310810725328,-0.00103583266932272,-0.014916033180699
"3057",-0.000715523978348842,0.0072548627968656,0.00345510773573321,-0.00344669189982472,0.00495013551740797,0.00296816771781572,-0.00272621893719094,0.00442825355766496,0.00167503385957479,0.0044163819462697
"3058",-0.000429574226390783,-0.00348520045234024,-0.00525552400874585,-0.00853129121145901,-0.0113290203140183,-0.00353225782499245,-0.00285221864222474,-0.00440873058078584,-0.00708711566989773,0.00502508265366841
"3059",-0.00186267741809276,0.000932669974680334,-0.00965569345432249,-0.0130232705425546,-0.0034045593929749,-0.00258675562132749,0.00297966872268973,-0.00468894898846839,-0.00561395451737989,-0.00250004222829769
"3060",0.00624395897261776,0.00628936159265892,0.00294334278971964,0.00117815058745752,-0.00924299150729369,-0.00328135922452311,-0.00213896324450658,0.00209386033736414,-0.0170175097510687,-0.0112781954887218
"3061",-0.00363730176204591,-0.00416667744046073,-0.00311812637531717,0.00141214163180248,0.00783748657555861,0.00308939695420585,0.00416810677404356,-0.0036563645537615,-0.002625525171288,0.00316865365604024
"3062",-0.00136023824523646,0.00209199440237229,0.000919956730150995,0.00987085546988054,0.00209048498167141,0.000577650453076339,0.00308342365813674,0.00550471807957464,0.00131624714241929,0.00505365229360066
"3063",-0.00605686514777415,-0.00185572285264657,-0.00588235718694274,-0.0055854678535141,0.00367161167201457,0.00278983613921513,-0.00484743873642257,-0.0059960879155726,-0.000903713433259012,-0.00565681936947671
"3064",-0.00836557355215095,-0.0146408278947455,-0.011834347225558,-0.0184881508067788,0.00648462644032333,0.00335746978657459,-0.00178213213052392,-0.00131101082692786,-0.000822292567862037,-0.00252848771387459
"3065",-0.00200001665211735,0.000707486829128356,-0.00168413542342893,-0.00715302769837645,0.00421298163087092,0.00143438717559063,0.000952072043749252,0.00709020871740162,0.0109455516262769,-0.000633692099297978
"3066",0.0145013686052557,0.0084845599938248,0.0108716157044206,0.0187319268412474,-0.00296131002422406,-0.000763802764126686,0.0147444263906507,0.00547598081210521,-0.00488438635247102,0.00126825226655392
"3067",0.00377101549159442,-0.0009348495331849,0.00241062258063818,0.00518625724912858,0.0070125958199776,0.00277083144336654,0.00410128198102999,0.00233390535211297,0.00605370592365362,0.00633316485474422
"3068",0.00661936286871589,0.0109941935053683,0.00388443427664797,0.00117259997660124,-0.00188431031468506,-0.000381053958764976,0.00455125776710608,0.00569230206449967,0.00699294990259514,0.00629318041424543
"3069",-0.000640074176765149,0.00439613657079652,-0.0106872603304083,-0.00538763254386698,-0.0072230826529941,-0.00142978618971712,0.00151013434222214,0,-0.011547093396224,-0.00437765136383261
"3070",0.00494080799075158,0.011057242989378,0.0115477973333267,0.014602036991525,0.00661433738231287,0.00315000993573533,-0.00231984587186362,0.0051451598173502,0.0045747649840775,0
"3071",0.00362581459646494,0.00455702704076466,0.00276186484599905,0.0111419754015512,-0.0005750245422802,-0.00133223494706203,-0.00558070965224977,0.00295659729088626,0.000569244526557489,0.00502508265366841
"3072",0.000247868158327114,0.00362887825024916,0.000367303963107135,0.000459119317771206,-0.00221870703506355,-0.000666966893372978,-0.00292279647891269,0.00179464181546396,0.0027632964664881,0.00250010572949733
"3073",-0.00300988684759818,0.000225929747827314,0.000550592436893149,0.00160631217137341,0.0104603054872079,0.00696044959436204,0.00334202276287643,0.00614111947671647,0.00648405754135339,0.00748116896669782
"3074",0.0112947147179681,-0.00271123505062421,0.00660430747930185,0.00137451796693067,0.00220068047901534,-0.000473608424877092,0.0169491102171229,-0.000762897674842389,-0.00402641327105813,-0.00495051590324702
"3075",-0.0192463230141504,-0.022881692576062,-0.0107527035612419,-0.0292839008386429,0.0155349010062411,0.0073892986424644,-0.00601852885186671,-0.0106897177419757,0.00234476875808531,-0.00870642553817436
"3076",-0.000752039209287791,-0.000463788846530644,0.000552754440652947,0.00235683169886514,0.00160192849313567,0.00253894276458899,0.000232921785329188,0.00643159858090558,0.00766312004788983,0.00376411527292286
"3077",0.00745415678964245,0.00417547419614883,0.0110477067180161,0.00305661074142627,-0.000719869943612617,-0.000844142019053584,0.00745070469557985,0.00409001782908147,-0.00496313648676172,0.0018750634218232
"3078",-0.00522924565794503,0.00207894651065832,-0.00346021711902722,-0.010782867252812,0.00920238811391938,0.00291016726045967,-0.00208016178296133,0.00127290472138508,-0.00522929190918853,-0.00561453565263736
"3079",0.00379044535391881,-0.00437992210146476,0.000548253088611395,0.00663494177477819,0.00348847585184364,0.0000936977245378223,0.00868461946934951,0,-0.014152850559598,-0.00313672023395206
"3080",0.00630565316533804,0.00463066489889985,-0.000547952671866692,0.010357938468734,-0.000947936125162196,-0.00159125887041123,-0.000803636378882033,-0.00127128649480368,0.000902378984374508,0.00062924131247688
"3081",0.011859173960961,0.0124453698425624,0.0126096133235207,0.0165423458615164,-0.0142042004383038,-0.00687637374620242,-0.000344647555551414,0.00305498271585858,-0.00393412828564654,0.00943396226415083
"3082",0.000489781696696667,0.00318684839665795,-0.00685791243329958,-0.00320867902600519,0.00184943596148446,0.00170264758778393,0.00643605556595594,-0.00456851733230046,0.00370282237885977,0.00249225404025921
"3083",0.00157360764362169,0.00816881960973892,0.00599673558421809,0.00689816240179364,-0.00866774185432218,-0.00311623414107942,-0.00102775721945936,0.00382452763573315,-0.00147565170989539,0.00124302907589291
"3084",0.00265339316190172,-0.00135056099085473,-0.000541896223168248,0.00616580621478957,0.00283345691861014,0.00104196264472534,-0.0014861499820451,-0.00482591820981704,0.00254513951038238,0.000620774470232011
"3085",0.00484018296027044,0.0015777299674431,0.000722926270185553,0.00771666824789929,0.00129161932867317,0.000473298530137445,0.00686892392795668,-0.00765703530851225,-0.00106459748534438,0.00310163159940502
"3086",0.000762501984449271,0.00180018475630317,-0.00234778042478234,0,-0.00354733178116295,-0.00160801699462243,-0.00591237678967915,0.00282940808552823,0.00434496628107151,0.00371063797274185
"3087",-0.0051248681128141,-0.00539087341361766,-0.00543099558201321,-0.00202698496309517,0.00315557804571931,0.00180001513321915,-0.00480383224853209,-0.00641211868611491,0.00522406325648417,-0.00184842871977575
"3088",0.00341101950573885,0.00338760240092939,0.000182094467796379,0.00473930875171646,0.00241970902515831,0.00236429519526715,0.00907936555998834,0.00877660204586905,0.00308564347404561,0.00864193295515259
"3089",-0.000277643727650378,0.000225038156040025,-0.00309380129171399,-0.0107817526495073,-0.00587398832326425,-0.00226425745666892,-0.00102506498233457,-0.00332662089414981,-0.012790431577677,-0.00489591927758426
"3090",0.00676593771993206,0.0063006940727619,0.00511136791719857,0.00726612973107321,-0.00712247744963912,-0.00463338968935589,0.00524471741665122,-0.000513401097571031,-0.000983968863894291,0.00307492641515528
"3091",-0.000654850630425918,0.000894433115869342,-0.000181622535562087,-0.00518480680281652,0.00252718879560576,0.00133028040313454,-0.00510381602099008,-0.00411000772234626,-0.00188790935093308,-0.0018393001365179
"3092",0.000655279740777281,0.00022335548257546,0.00399644039253899,0.00747789331392568,-0.00626116927927434,-0.00341531853275989,-0.0214321024056161,0.000773749128404111,-0.00896378304216749,-0.00368550360883424
"3093",-0.00244691782599005,0.00402056012163898,0,0.00292399442219327,0.000409007486621205,0.000190259380052238,-0.00908649968923747,-0.00541231564587974,-0.00190858016913809,-0.00369913679082623
"3094",0.00196926367188599,-0.00200219480911934,0.0014473847597003,-0.000672899907299684,0.00523482492269478,0.00237951844528173,0.00681876959238159,0.00155480333384772,0.00074828733578558,0.00309401742611271
"3095",0.00086177792826736,0.00044580914736092,-0.00361330683492844,-0.00650807767785277,-0.00480071868797893,-0.00142442709001123,-0.00980856465799673,-0.00155238967320848,0,0.00493537152270385
"3096",0.0089917074152055,-0.000445610490128256,0.00562103506005718,0.00225887454993323,0.00212601314788685,0.00180631922048735,0.0119103338370743,0,-0.00207692941571169,0.00122758060901673
"3097",-0.00221917283369477,-0.00557296670460128,-0.0122611813086461,-0.0135225597912375,0.00815831151980118,0.00379693456129915,0.0065261588757286,0.00207310973877184,0.00291373619096569,-0.00367860027303579
"3098",-0.000615895766010288,-0.00201743122183107,0.00219064822687787,-0.00137084516990382,-0.00145671111425838,-0.0012292957592881,-0.00196837686737927,-0.000775836727594847,0.000830073870423442,-0.00184621621650349
"3099",0.00465667126144975,0.00134773610608407,0.00910742283635302,0.00388937313179993,0.00340392329672179,0.00265060886085577,0.00754072384556959,0.00258794715121846,0.00663517458737672,-0.01171384965108
"3100",0.00156767248773559,0.00471056208501497,0.00397111747043821,0.00205102948781533,-0.00638070485466968,-0.00207709970974812,-0.00955674460749478,-0.00154878326768071,-0.00444921303989754,0.00062387250715612
"3101",0.000510506504268537,0.00468857083453433,-0.00359582227192756,-0.000909866685288696,0.00512127034984311,0.00198690821747327,0.011392689977324,-0.00258515538187665,0.00306211200757911,0.00311710095042761
"3102",-0.00751650887797395,-0.00755559896687419,-0.00342830019713147,-0.00751181970794712,0.00412502043691276,-0.000454195856966377,-0.000689696950093799,-0.0028513223888863,-0.00660061897526276,-0.0031074148247241
"3103",-0.00215911325323503,-0.004254295181219,0.000362052125365775,0.00229358634399479,-0.00476188742722994,-0.0028397934920894,0.000345128973241682,-0.0122172498247209,-0.00382059794317935,-0.0112220701642258
"3104",0.00978794057695564,0.00966950093668917,0.0128506299927442,0.011899361572911,0.00283844979489589,0.00132919449269964,0.00793368634698099,0.0202630750850943,0.0059196263811967,0.000630495656581909
"3105",-0.00411519042438591,-0.00913139127331453,-0.0101858021289634,-0.0205789998100873,0.00274929148837644,0.00255951183209535,-0.00330811788605612,-0.00412696959926884,0.00132611684498762,0.00315068397557128
"3106",-0.0166998115375983,-0.0188807427840351,-0.0182343078420995,-0.0196259640551943,0.00766129774970015,0.00340433147114871,-0.0181984743293513,-0.00207192020842906,0.00331099252232425,-0.0125628342747678
"3107",-0.00138917938247973,0.00504005667773288,-0.00606841428840321,-0.00141304076352511,-0.00432179782543618,-0.00188502863681028,-0.000116602804605015,-0.0028551098763212,-0.00247500208295515,0.00127222146063866
"3108",-0.00302572424128678,-0.00569863434887896,-0.0064754975809459,-0.0158018626911457,0.00409938765774487,0.00264399514517066,0.00233178656205424,-0.00025996531526129,0.00239842023328363,-0.00508254897919436
"3109",0.00502344891777273,0.00664845283713911,0.00689014751737305,0.00599072745460605,-0.00136077659978961,-0.000659089363468035,0.0105850231429283,0.00702924211873102,0.00189771456842536,0.00191564380807363
"3110",-0.0251302870659297,-0.021407478478418,-0.0225633268098948,-0.0333491153182287,0.00785568311663609,0.00499429468851531,-0.00115086401243003,-0.00646319193435452,0.010211628098493,-0.00509874586703907
"3111",0.00904368676772016,0.00791241946665244,0.0140019265445315,0.0140462946698072,-0.00294284531553934,-0.000937780405597666,0.00414836819340558,0.00468371328109929,-0.00171190187840398,0.0134529142144599
"3112",0.00585742429713854,0.00600324850424894,0.0014927397096276,0.00194403278739452,0.00614233825288335,0.00319089265414219,0.00654112780987859,0.000518153783467978,-0.000571615225964495,0.00884951432741188
"3113",0.00926125791062038,0.00895105220521208,0.00409914180511639,-0.00485077896938058,-0.00332991732176502,-0.00196446343352408,0.0059286508841927,0.0056947718951228,-0.00719010545951559,0.00563909774436078
"3114",-0.00646518847467159,-0.00636934811806844,-0.00371127600302401,-0.0180354569815251,0.00222723893965027,0.000468422391648016,-0.00283348962287222,-0.00669220069517351,-0.00707760666484059,-0.00934579439252337
"3115",-0.00661196336526815,-0.00663922366081937,-0.00540131737063521,-0.00421949449285297,-0.00206352347352345,-0.00168630633858324,-0.0147760329162724,0.00492346180819681,-0.0000829092402335752,0.00440255832365777
"3116",0.00901557356560456,0.00691402959249565,0.00692885580457836,0.0127118615349555,-0.00159071258808363,-0.00112616405109589,0.00842178570517449,0.00361013869264415,-0.00232093834815106,0.000626152843005601
"3117",-0.0030715011208382,-0.0038910247744095,-0.00818301676629962,-0.00492259212176771,0.00573566289970961,0.00300649635178174,0.00354653247096137,-0.00693724853411204,-0.000997033890021259,-0.0143929485468923
"3118",-0.0122185152161854,-0.0101101270890894,-0.00750047392013242,-0.0128616868452219,0.0112475317072567,0.00608930756106707,0.00136796352520818,-0.000776122523459155,0.00773453106677535,-0.0209523796007606
"3119",0.00226843799230059,0.0106776149556274,0.0154921750349151,0.0010023217177566,0.000861637101620794,-0.000279634552242891,0.00330135060189596,0.00828576522543956,0.00107291410535471,0.0136186761454711
"3120",-0.00930057573396836,-0.010564808003684,-0.00837216836311616,0.00350435147966022,0.00719997219398461,0.00437766173973397,-0.0105525678785896,-0.0118130951388754,-0.00387469899732817,0.00831731624288978
"3121",-0.00671057023511235,-0.00928529416045465,-0.00469045685272296,0.00648539535182224,0.00303023589319551,-0.000371014617387089,-0.0119264568168406,-0.000779580448413975,0.000331051885607003,-0.00380710643535986
"3122",0.00273110209572458,0.00585762215305086,0.00452405692150615,0.00545239566003142,0.00859855973831225,0.00361775190674152,0.00406214303863828,-0.00182054683686317,0.00678413981672543,-0.0101910607913405
"3123",-0.013475236725235,-0.00931756727499489,-0.0106961429716511,0.00345071963417243,0.0125193283948097,0.00665502210306124,0.00416130325942832,0.000260556628771891,0.013476867228583,-0.0263835464521808
"3124",-0.00254296313024627,0.00705401215013346,0.0058801230950245,0.00908880488409514,0.00668844404001523,0.00481140363290611,0.00391398565698586,0.00859615809224268,0.0144328141663372,-0.0033047148998443
"3125",0.0217066793987741,0.0121408567314394,0.0115028846939802,0.00219072516638441,-0.0114010420343447,-0.00366211244096915,-0.00321078680676734,0.00413206723473247,0.000319726638000839,0.00596816962723756
"3126",0.00866208968617466,0,0.000559272491531537,-0.00801553190458137,-0.00565179566963436,0,0.0209365260446996,-0.00411506351561075,0.00255692365070836,-0.0204350464341544
"3127",0.00650260575430583,0.005536468731421,0.00111795826643379,0.000489799722949602,0.00322590690151259,-0.000183946760951681,0.00146470490990236,0.00335708808101054,0.00326768149145074,0.0174966572558402
"3128",0.0100070939339316,0.0126175207104506,0.0120975359921032,0.00783155124848167,0.00865180855606096,0.0039522528201803,0.0030377443875933,0.00566310063342224,0.00564028453225962,0.00330683328664261
"3129",0.0045888827531213,0.00203893646701747,0.00459728412761473,0.0104419574489978,-0.00941239408945627,-0.00494362601179521,-0.00302854444370693,0.000255955010062703,-0.00995334576043438,-0.00263676074053543
"3130",-0.000242176198560373,0.00520009233786545,0.0032949000205087,0.0112953958561104,0.000613049425299605,0,0.00168762257545807,0.00511761863525617,-0.00119685628027033,0.00660936264706513
"3131",-0.00176527864315279,-0.00584789763405991,-0.0111293002776259,-0.0106938684862097,0.00076565537408535,0.00257606868498406,0.00325730717078132,-0.00865583179715668,0.00519253874420822,-0.0137885081622434
"3132",0.0041262316787587,0.000905027410576631,-0.00110715954658069,-0.00168157872299102,0.00344341082415967,0.0024776356475269,0.0036945631326637,0.00308165702068619,0.0061193355142759,0.0126497765772546
"3133",-0.00110486058397807,-0.00791154357945911,-0.00258580940943687,-0.0110683407622449,0.00251681031126094,0.000732443700612428,0.00167321021861522,-0.00409632910581226,-0.000315955771184151,0.00394477291203388
"3134",0.000380286135369445,-0.000467642879882102,0.00293384177610134,0.0039471732586942,0.0017493598832774,-0.000183030663175598,0.0107166486057249,0.000514175993955979,-0.000632071754615549,-0.00458419598484128
"3135",0.0104709263228921,0.0142722191536424,0.00596237888521411,0.0241758178254665,0.00501209853753148,0.00192139297310945,-0.00177639610018565,0.00668047936755345,0.00506008843152861,0.0118421049993025
"3136",0.00225722138052675,0.00438305478385059,0.0088906068585628,0.00834530573057068,0.00143535978788556,0.00273949262445505,0.00622841559506315,0.00280754347008538,0.00605723711318662,-0.00195051907153276
"3137",0.00955425752788464,0.0101056269928825,0.00973010836657839,0.0146606571605734,0.0026406384642268,0.00163914355486883,0.0044214015220152,0.00763562648919791,0.0251779030821637,0.0201954158937032
"3138",-0.00145353266300652,-0.00159168521422848,-0.00981829524999533,-0.00326267209768072,-0.0109865530756981,-0.00409119471570296,-0.0126555423018347,-0.00303106101932626,0.00663561126812895,0.00255425662399422
"3139",-0.00122442405360756,0.00159422271495191,0,-0.00140281312967272,0.00745671943877224,0.00346882527491643,-0.00624160607219082,-0.000282025293394716,0.0148507808713678,0.00445857696222429
"3140",-0.00980816784632088,-0.00568441997332425,-0.00440676127949446,-0.0103020879290587,0.00309655404383835,0.00154670622955688,-0.0127861382476872,0.00102514813054744,0.00194113032789112,0.00317059845271306
"3141",-0.000997256938596203,0,-0.00147557334342474,0.00946290730533406,-0.00639995976707464,-0.00408769207058213,-0.0188592879495546,-0.00512040648066303,-0.00916539513782555,0.0050568469803165
"3142",0.00354590776452812,0.000228717074466589,0.00406363875874938,0.00703089332949447,0.00704728711792901,0.00300998497361316,0.0115795210919611,-0.00257332309398028,-0.000977701729880986,0
"3143",0.00514578181644776,0.00754455272130206,0.00404709824688854,-0.00139640447827205,-0.000677253872796602,0.000454728022696527,-0.000572383304704771,-0.000257870718607278,0.00271003470972686,-0.0106917812989837
"3144",0.00907861187880177,0.00294989353359587,0.0142909198828265,0.0118852859506371,-0.00233868426474104,-0.00125654568743028,0.00343608673166784,0.00335475316468092,-0.0193693848206319,-0.000635706350688436
"3145",0.00260430701466841,0.00316733966440452,0.00307077176439252,-0.00253333572691083,0.00771310409689785,0.00355553467891556,0.0156375113469689,0.00488692362148435,0.0213597389894249,-0.0165393960464058
"3146",0.00799506493414937,0.00721693762029751,0.00288137929147259,-0.00184716850054689,0.00712923050620118,0.00190770214372971,0.013261436253716,0.0133095578577602,0.00164905924146463,0.00970239117406657
"3147",-0.00113784955242147,-0.0107478054572476,-0.00430957764988016,-0.00693964665337143,-0.013263157455524,-0.00634713350804106,-0.00454749709149749,0.00176783738934194,-0.0111502353083054,0.00192190997549258
"3148",-0.0054947775173072,-0.00452693563301965,-0.00577098014921029,-0.00605644282582773,0.00135936475824283,-0.00100350223097889,0.00323101388653213,-0.00352999281323829,-0.00643261697012709,-0.00127885885720846
"3149",0.00124641666598935,-0.00409282813497358,-0.00888807915921874,-0.00304653963394874,-0.000377056924528052,-0.000639407479482212,0.00488692721289685,-0.00328939031474451,0.00350374761616434,0.00320104594039505
"3150",0.00477818322040569,0.00365299199018598,0.00603947320362197,0.00846260555322442,-0.00550661086927295,0.0005484008921679,0.00530494692702965,0.0020310933994796,0.0157874914611007,0.0216975534556096
"3151",0.00234409463059659,-0.00159240942167171,0.00181918487105803,-0.00186474957494176,-0.0133511820766316,-0.00493285622037376,-0.0112136459804788,-0.000253540108381523,-0.00844358501914999,0.000624588412292182
"3152",0.00447705796967646,-0.000455602872050043,0.000363157695488336,0.000700502674902292,0.00115326061263565,0.00110162546680459,-0.00177905687298552,0.000760420992281352,0.00625472508488456,0.00249679418045523
"3153",0.000332375148266895,0.00182356979760079,0.000726144655517125,0.00373394803941807,0.00575975518701233,0.00210902476751684,0,-0.00202597789148029,0,-0.0105851998891362
"3154",-0.00322496947150397,-0.00341302214203532,-0.00743693652346356,-0.00139500951081428,-0.0029778592083195,-0.00219625997290185,-0.00233899574470953,-0.00304484167050523,-0.00846255529440998,-0.0106985729502709
"3155",-0.00680519656894341,-0.00205478894955691,-0.000913785450541549,-0.00302667850066507,0.0107979744800613,0.0046773192161591,-0.0040193666164352,0,0.0164653179667065,-0.00890587338578497
"3156",0.00366097461390136,0.00503320909893112,-0.00256081579297918,0.0060720250548234,0.000075645959967563,0.00246448268685961,0.000224407373496494,0.00432672091898789,0.014117951937614,-0.00706035519196246
"3157",-0.00555497595686383,-0.00614619478306921,0.00256739040687992,-0.00510685096893992,-0.00234831276814973,-0.00182085657648656,-0.014681274854097,-0.00405470077845793,-0.0147273963870866,0.00581777724944499
"3158",0.00245641895389981,0.00206144839882971,0.00146333401310583,0.000233250678514318,0.0018984477532471,0.000455960769112806,-0.00181983634482952,-0.00559787626312769,-0.000148761804500963,-0.00321338909511093
"3159",0.00715019139277406,0.00640002402989293,0.00803648336285101,0.00116636879585785,-0.00545717000028323,-0.00164128374433958,0.0101414175065579,0.000511490024671657,-0.0056526219186156,0.0064474309978213
"3160",0.00469947561725936,-0.000681429447965343,0.00126831611461853,0.00163095591273033,0.00434360905644193,0.00146126555097825,0.00281991635238721,0.0015347317601031,0.00508634146029863,-0.00448428304224902
"3161",-0.00477692665449392,-0.0104544652514237,-0.010676734376145,-0.00883930614960748,-0.00477993314794156,-0.00173280810958587,-0.00461195053674535,-0.00561803018370721,-0.00707000844943095,-0.00386106898946703
"3162",0.00669977483057527,0.00528250505800121,0.00256079706302303,0.00211215748171378,0.00236353157130464,-0.000182691957795633,0.00339036202044518,0.000513584552739532,0.00164893571651836,0.00129201154218861
"3163",-0.00182118337756088,0.00182775944459257,-0.00127709070148163,-0.00187348374662444,0.000304022442131568,0.000913691960279017,0.00292825176214784,-0.00359333156116071,0.00665968277955487,0.00387103320698201
"3164",-0.00245456715467229,-0.0150514170882696,-0.00639388062250812,-0.00774285748866399,0.00243381898215023,0.000456359088098823,0.00718698535199147,-0.00644004998621805,0.00334495654013933,0.00578399589622292
"3165",-0.0109404657117587,-0.0064829117450278,-0.000735471279400324,-0.0122961229163161,0.00804004118390189,0.00255528676969896,-0.0033448252528514,-0.0111484238000432,-0.0131129726807816,-0.00638968965774234
"3166",-0.00870787101838777,-0.00419479076769436,-0.00018399372876432,-0.0196312861549998,0.0198607087560665,0.0113421126684405,-0.00100693237729022,-0.000524444055387652,0.0240221967708476,-0.0276527736668752
"3167",-0.00752947240716961,-0.0100633859799476,-0.00515264057731069,-0.00976801462671417,0.00924124096223267,0.00207380238217714,0.00447923668418682,0.00996838953012724,-0.0038120737830929,0.00132277363287803
"3168",-0.0300732039734811,-0.0217492198294577,-0.0247873228309007,-0.0369913296715889,0.0172880999165694,0.00863687814368341,-0.0179487929246326,-0.0199999597990181,0.0139818530722045,-0.00858656973011873
"3169",0.0140229948205639,0.00410818438029503,0.012708607477171,0.0143406912952577,0.00799317080018813,0.00160570728053488,0.0105574845709979,0.00477087770665485,0.00812839144276589,-0.00532973477973142
"3170",0.00059072143230221,0.00505412133123162,0.00693012012995853,0.0045442575372745,0.000357050887780597,0,0.0104470002710237,0.00501184788790998,0.0151896907295461,-0.0127260991363837
"3171",0.0196200343062054,0.0107758820972288,0.00706843711075678,0.0123146315413143,0.00214277604572621,0.0000891314803437293,0.0167871040165464,0.00524922129272531,0.00503468997206946,0.00542736221015194
"3172",-0.00681157546440514,-0.00497509460983592,-0.0105282091116399,-0.0101787847037084,-0.00199572442820029,-0.00151380321972949,-0.000109225769447829,-0.00365525316394311,-0.0033161716874669,0.00877197552943043
"3173",-0.012173077872124,-0.00785718640322242,-0.00952023346364483,-0.0120391796392081,0.0208499912324025,0.00633187849080197,-0.00382723683607544,-0.00445496034052772,0.00969849956457947,-0.00735781389097367
"3174",0.015551429300382,0.00863935935532667,0.0113079617057301,0.0126935902348058,-0.00342756387120702,-0.00354479467123148,0.00109759718901792,0.0023691566436157,-0.00595951742412126,0.0235847893992234
"3175",-0.0295675037760563,-0.0271235223513492,-0.024226620351416,-0.0288291617813374,0.0225295029915702,0.00667018181924584,-0.016227969601802,-0.0168067648948103,0.00684159265652129,-0.0151414293457932
"3176",0.00264176536135619,-0.000244426786795593,0.00954925205452373,0.0067112739993973,0.0111196931596225,0.00636093292387185,0.0110343385527971,0.00988250618086628,0.00665497022767081,-0.00802138964796029
"3177",0.0147548969052107,0.0119861946345963,0.0104048848829736,0.0138461916366319,-0.00801052440288685,-0.00263364527528032,0.00870910515329104,0.0134885086323775,-0.00640221307729039,-0.000673900029193431
"3178",0.0120478420110637,0.00773497527385869,-0.000187231950459443,0.00404652660358407,-0.014302316261108,-0.00475317982505674,0.00754103247567661,0.00287050372352216,-0.0116963020849999,0.00472013878150723
"3179",-0.00766261728266371,-0.00575665424371397,-0.00205999466731954,0.00201516139670233,0.0103447898982616,0.00442217424071245,-0.0074845909323884,0.00286220121468705,0.00779537943593356,0.00268454096763349
"3180",0.00813550104661487,0.011821367336702,0.00337784126751584,0.00955237490071648,-0.00666553262411473,-0.00264152956252139,0.00371579558562307,0.00337326291847306,-0.00316441866147987,0.00334674288307091
"3181",-0.000307781162403042,-0.0021459170209025,-0.0014962513858594,-0.0129481814042265,-0.00664090417500462,-0.0022072186613542,0.00555323612958403,-0.0036203931307186,-0.00253951052975143,-0.00466975715446305
"3182",-0.0256875819349763,-0.0126641261072956,-0.0112379916934224,-0.0148838404967545,0.0164346432924856,0.00672458018323652,-0.0137520725807214,-0.00207631314454215,0.0195898452442651,-0.00737260842225429
"3183",0.0110585966816674,0.00701838699270629,0.0145860646303937,0.00537766288708008,-0.00404252453587428,-0.000966819133274455,0.00735609868994436,0.00520152547181318,0.000138752863130476,-0.000675265120282376
"3184",-0.00392351092850196,0.000480666040632016,-0.00317404820279221,0.00178310710113516,0.0154090624328171,0.00431084492386669,-0.00381472281823769,-0.00051732366381041,0.0095707398630871,0.00675673356420781
"3185",0.00704143297489668,-0.000720714322002269,-0.000374604198213668,0.00279667611022494,0.00128730267190313,0.000350204033951806,0.00229763048096632,0.00232981963944945,-0.00281653486490541,0.00872487747592454
"3186",0.0127728514278389,0.0100960931440408,0.00712016618920552,0.0111563219030255,-0.00378909358803536,-0.00192646458053713,0.00796858863462235,0.0005163597825939,-0.00716456993208681,0.00266132126566654
"3187",-0.000444197610582897,0.00356971094291092,0.00316269489205223,0.00777324461046813,0.000271560777266533,0.000263215303470066,0.00129947714861123,0.00438829118585726,-0.00256727041934735,-0.0159256794434508
"3188",-0.00584722669212823,-0.00308263298410483,0.000556440100536459,-0.00622039468323821,0.00129251550097398,0.00219657308406673,0.00973402501557707,-0.00565423990284786,0.0139130434782608,-0.0053944247471307
"3189",0.011350445959456,0.0164129591746451,0.00556073707382021,0.0167750942965141,0.00149462118021293,0.00157779566429705,0.00781905163935526,0.0129234080646554,0.00624359519725548,0.0237287654582146
"3190",0.0128552604024939,0.00514854762317052,0.00718892553148121,0.0113272485527247,-0.0181101475791023,-0.0080524336236325,-0.00627047890575572,0,-0.0240011243965328,-0.00132452568052432
"3191",0.000772444040410214,0.00209543014511748,0.00347732639974452,0.00438278999241848,0.00711491216826787,0.000617622156134257,0.00192508337356312,-0.000765547010674106,-0.00852313125976756,0.00265256475118081
"3192",0.000503225849771693,0.000464624435777106,0.00656567500515681,0.00315161548600229,-0.0177650421605977,-0.00617282179493883,-0.00651144260716663,-0.00229817471751481,-0.00373449131531134,0.00925928103607609
"3193",-0.00023480660068198,0.00139348825050623,0.00289905597094231,0.000724779396400033,-0.0175281322829872,-0.00727593001834015,-0.0106371746751081,-0.00307145166505018,-0.00855793202176902,0.00131050490558815
"3194",0.00711109353226891,0.00533386298470706,0.00885282626573347,0.00700323195049002,-0.00177677720061453,-0.000983199132127299,0.000977254564115126,-0.000256839854801516,0.00606367557744147,-0.00719890871020412
"3195",0.00346385424453866,0.0059977771870654,0.00662605836786168,0.00719434165689492,-0.00655087967380963,-0.00223678813089701,0.00488254789522791,-0.00154078204874075,0.00205635681809802,-0.00395517459858208
"3196",-0.000663857007232149,0.00275166273805172,0.0117416609789243,0.00571419915139715,-0.02135890855775,-0.00914619525039095,-0.0116606720238926,0.00823057378409597,-0.00827917451207039,0
"3197",-0.00308884500471585,-0.0107477538736637,-0.00527509414390059,-0.00781248982579141,0.0127438232539892,0.00434386678732457,0.0102687984435916,-0.00433676714081166,0.0083482914740618,0.0443414722905136
"3198",0.00253201543524373,0.00485433966964077,0.00371209171729014,0,0.00542320602547108,0.00261283430491921,0.0109210677808038,0.00614908562765315,0.00198131181807826,-0.0190114068441065
"3199",0.000598133530704814,-0.000920127700753892,-0.00211341472372228,-0.004056234525186,0.00424370761096138,0.000359669801191398,-0.00352950147708941,0.00050926866148715,-0.00628530340599009,-0.00645992644230764
"3200",-0.0000665000076969235,0.00345388716909478,0.00741273493675521,-0.00407282917093665,0.0030083623973669,0.000449379933336713,0.00483022178791992,0.00610839464331847,0.00405082774247889,0.00520164843502324
"3201",-0.00472478623974903,-0.00206523231749223,-0.00227750059499665,0.000962155379854446,0.0132103373071777,0.00574700506325354,-0.00042728243259138,-0.000758962528595308,0.0118204842286274,0.0012935513870731
"3202",-0.000234707890673813,-0.00252925235923485,-0.0010536517886981,0.00096140513265075,-0.00021130637677591,0.00142853916137908,0.00149616696422239,0.00104781563549827,0.00559638346826974,0.00258408871869475
"3203",-0.00784659486491712,-0.00576304225355295,0.00140624886099672,-0.010564252297264,0.0120541182253315,0.00499286350446471,-0.00124662170224565,-0.00357407606328586,0.00528692173913048,-0.0115980023440451
"3204",0.00591461935143722,-0.00486906630152562,0.00403729029037625,-0.000728071511391426,-0.0146270936510212,-0.00656489536216209,0.000753197564228092,0.00358689590207084,-0.0185453815841596,-0.00586701408252943
"3205",-0.00208317900438204,0.00535881357581092,0.00174819031350837,-0.000242842124415721,0.00643277259655806,0.00214322775649833,0.00817218092955807,0.00638239051935185,-0.000282091232008841,0
"3206",-0.00538722028828265,0.000463439979490499,-0.0143105868989339,-0.0128734815718351,0.00245792589385507,0.00142567518426095,-0.0060794505316254,-0.00329770968614373,-0.00514842397939885,-0.0039344926789654
"3207",0.00463771776021304,0.0023165545873729,0.00460331744523157,0.00565945641023347,0.00245223577403841,0.000800938021435549,0.0037557263283674,0.00585379047943335,-0.0155253298670827,-0.00987485104181107
"3208",-0.0118947351094091,-0.0108620826985468,-0.0044059985103938,-0.00709555941158391,0.00301046870471255,0.00276947939558791,-0.0105837204102077,-0.00657903542414928,0.00547281650006548,-0.000664871068921102
"3209",-0.0176645744498442,-0.0261682261822015,-0.0123916460562183,-0.00763936170484869,0.00244302436427057,0.00346320820901691,-0.00388963676821408,-0.0056035309257545,0.0116736370524373,-0.0086494124123877
"3210",0.00819258813739276,0.00695784176502712,0.00501886859219636,0.0129128121322655,0.00912206246348357,0.00522109577092866,0.00976228843180804,0.00768443375981476,0.0045306457783747,-0.00134230457842133
"3211",0.0135322410685474,0.00905397622871673,0.0115926834759006,0.00441300283682855,0.00738343920600615,0.00193691689071107,0.00537114787806559,0.0119471679895657,0,0.00806451612903225
"3212",-0.00431473988080566,0.0002361942027862,-0.00634702262289311,-0.00829880059754284,-0.00828806387283121,-0.00333883554191061,-0.00277805455035196,-0.00326540326940861,-0.00852707576576783,-0.0013333559115386
"3213",-0.0155246621108315,-0.0110953311169494,-0.00585523276420208,-0.00713754881971296,0.00269353889327117,0.00211582657828036,-0.00514307307233053,-0.00302425675985984,0.00874259707523506,-0.000667466324014487
"3214",0.00949650681304526,0.00811640985309836,0.00874529353149267,0.00768470873433569,-0.00564846398384988,-0.00255120461856251,0.00323099192944287,0.00505540397983828,0.000916044263191251,0.00267198788324197
"3215",0.0067633230526063,0.00899833107529635,-0.00123838016504674,0.0103319914667417,-0.0148946193035843,-0.00626228529716577,0.00193242543626693,0.00100617687383031,-0.00872935567625432,0.00666220231940717
"3216",0.0103669218286517,0.021121768414923,0.0124002992993675,0.0160702047005306,-0.0123766385660564,-0.0068340458457341,-0.000750047508989438,0.0100502516710979,-0.00553937228235746,0.0119126403683329
"3217",-0.00111378239557602,-0.00436684231472229,-0.00437446090573157,-0.00431347162050699,0.00726266505335604,0.00277035437837991,0.000214490413857904,-0.00124372325531197,0.00399912164535543,-0.0045781334059144
"3218",0.0099003186472022,0.0129271751210032,0.0149384142524358,0.00890484626842047,-0.0120879868634084,-0.00481234922362528,0.00053600512070906,0.00697381249166518,-0.00697058843361797,-0.0026280985247561
"3219",-0.00160591669150634,0.000911553673747401,-0.00207784576542747,0.00286266388577427,0.00121648992525092,0.0019700097942279,0.000749969502087167,0.00692559650910662,0.00573026999691795,0.00131747834751383
"3220",0.00294898607001959,0.0047814853839514,-0.00260286183318859,0.00380596522259435,-0.0024301403891982,-0.000357477711380838,0.00556748983340727,0.00147372229113985,0.00142437856493483,0.00394743517647012
"3221",-0.00437717595740506,0.00067969915030397,-0.00191372043456384,-0.00521341872605818,0,0.000893950331277926,0.00798559958052292,-0.000245218646040102,-0.00106673777777744,-0.000655352323614466
"3222",0.0067791037050291,0.0040760758059335,0.00714656325024943,0.009052071955723,-0.00752251416383287,-0.00366226920308088,0.0072884145956682,0.00588824938058319,-0.00477014072767334,-0.00131149755965509
"3223",-0.00326670272927365,-0.00405952885856964,0.00121151680138443,0.000708011628385519,0.00584707688677155,0.00233111480080717,-0.00325079319181554,-0.000731796062110823,0.00293299964611915,0.00131321984427624
"3224",0.0029097444658559,0.00634060369601785,0.0041487380295675,0.000236130717597316,0.0010049427050236,0.000357629234640333,0.00136768578837132,0.000244021558685859,0.00235379462953911,0.0124589936319914
"3225",0.00163400135241698,0.00360040657338145,0.000516425401974274,0,-0.0020075312257507,-0.000178891392962899,-0.00126086162348826,-0.00390432776182037,0.00711591835989411,0.00518143477574506
"3226",0.00409482762880775,-0.000672651525742252,-0.000516158844435566,0.00707539508593436,-0.0048850978845979,-0.00214614565428906,-0.0102041250618702,-0.00367473984778377,0.00233167527966982,0.00579890297429775
"3227",0.00563651971534029,0.00426282491603991,0.00292640473543959,0.00585474608954972,-0.00909624974703416,-0.00376410786393633,-0.00542032359649225,0.00122945804967856,-0.00860004223459732,-0.00384362468784738
"3228",-0.000296645385901684,-0.00134037960242139,0.00429109916276227,-0.00512218841846956,0.000655962963953094,0.000899499285002658,0.00341955583206399,-0.00122794833870898,-0.00277303045202659,-0.00192926024006812
"3229",0.00306726146369174,0.00626391370257884,0.00273460905837641,0.00444658217165461,0.0146337529295297,0.00485364997144133,0.00553785511493987,0.00442591972660566,0.00549022459893056,-0.00644334190948614
"3230",-0.00266334645185196,-0.003334798849566,0.00017051568148263,-0.00792173404246355,0.0134903779901219,0.00635043202688523,-0.00169440166600887,0.00342719556542281,0.00999850347472697,-0.0058365754909161
"3231",0.00926395994162621,0.0073611831390592,0.00988405287611704,0.0150304743322298,-0.00307807722415476,-0.00188700316004742,-0.000742658226989157,0.00390337517356243,0.000912764209712646,0.0182648168799422
"3232",0.00401764672577709,0.00465019580232462,0.00674997279386402,0.00994919104212344,-0.0131615709019579,-0.00508338862162339,-0.00775041220686645,-0.00121501033573157,-0.0028760101413583,0.00640612793002915
"3233",-0.00110612204278604,-0.00264498751151609,0.00134093979578842,0.00572741793487364,-0.0112465527501098,-0.00537826568941457,-0.0162635830741514,-0.0036496783116462,-0.0161800077177632,0.00254619201042838
"3234",0.000227922288821958,0.00132604638945666,-0.00217607485604265,-0.00318925997110975,0.0060516197653544,0.00288388839653564,0.00293656553507815,-0.00293027734405138,0.00429024650882015,-0.0107936716004128
"3235",0.00351680021171541,-0.000220854782100766,0.00587142919547223,0.00731276554429616,-0.0181184969415058,-0.00799781318243531,-0.00954324036171261,-0.00269424542875596,-0.0155214884055853,-0.000641891971205011
"3236",0.00246624008727125,0.000220903569710496,-0.000500251116052786,-0.00907450823603551,-0.00420727568287393,-0.00135883555657179,-0.00186137120989693,-0.00982318329241527,-0.00636439556333568,0.00256908653475652
"3237",-0.00190977160134997,-0.00154496383120561,-0.00250303712978517,-0.00709702522355227,0.000667268337769533,0.00108861564954355,0.0023036368681888,-0.00471229439952836,-0.00240192883326229,-0.00640612793002915
"3238",0.002107747975028,0.00110523371805682,0.0021746361072601,-0.00645601413047459,0.00459234727806024,0.000453003984913991,-0.00700445069906486,-0.00523302784300372,0.00269951120238598,0.000644788954934805
"3239",0.000323828465847331,-0.00198718807514875,-0.00350514194194318,-0.00765847513892637,0.00648866627475853,0.00271717880993871,0.00815590673709021,-0.00551099646610509,0.00400205943399845,0.00193298947981591
"3240",0.00145568995157896,-0.000221278697407623,-0.00435523711165187,0.000701558465661112,0.0103299086046611,0.00505811397596179,0.00798070152959029,0.00428214854773112,0.00420352237146027,-0.00321552085191401
"3241",0.00723649644061464,0.00464710867952078,0.00588837738977332,0.00794582603030336,-0.00108784040890453,-0.000808778748280892,0.00531463568713697,0.00777521560686112,-0.00252591660689849,0.00516131205968251
"3242",0.000737548232146334,0.00132157462605664,0.000836230890151279,-0.00162301487261485,0.00181500486757025,0.00170895986198705,0.00517850590718383,0.00746640862929393,0.00296641327859848,-0.0102695541958202
"3243",-0.000288456745617061,-0.00131983037172667,-0.00317510104484298,0.00209018080705148,0.00833267159737971,0.00188563174388734,0.00128797352944754,0.00370557784018444,0.000505028152684606,-0.00907920528324691
"3244",-0.00371863188994093,-0.00594718757947343,-0.00301756884768256,-0.00440342140464778,0.0103478194781796,0.00367461361614763,-0.000214421435213552,-0.000738352491468697,0.000504672283442753,0.0130890276901821
"3245",-0.00160901419779902,-0.00177267964951355,0.00100881461888958,-0.00209485315733615,-0.00625883871237065,-0.00250033172801323,-0.013723617875501,-0.00492601403191495,-0.00547704689669382,0.00904394952668475
"3246",0.00222388708620636,0.00244173734341957,0.000671968496845254,0,0.0012881418482058,-0.000179167888932796,-0.00326111891551184,-0.00371294214239082,-0.00188402173913049,-0.000640183169661301
"3247",0.00775020580077079,0.00819301809070039,0.00688269951794318,0.0100302486958974,0.00293067959896787,0.00044767324725048,0.00392630059572152,0.00546592143956204,-0.00479165802266368,0
"3248",0.00226568905956626,0.00109828431465941,-0.00166730042884711,-0.00300221349964402,0.00584412277316071,0.00187945160670666,0.0120587717177538,0.004200457373154,0.00481472855537302,0.00576553466334007
"3249",0.00445757488852583,0.00153581206547249,0.00200401987316301,0.00115816718960327,-0.00290502239490109,-0.00259040910067465,0.00322007231439159,0.00196853645427653,-0.00529991268694952,-0.00509556275296941
"3250",-0.00370877100652445,-0.00569558805692871,-0.00949995369963796,-0.0157334240505786,-0.00213212673525776,-0.000806026426351303,-0.00278182970005747,-0.00294690926710228,0.00620397073950696,-0.0198463287199427
"3251",-0.0084947561324431,-0.00793121782771167,-0.00201919405982853,-0.000235102874464488,-0.0133329118892367,-0.00359037109241955,-0.0148068426320332,-0.00270929288186772,-0.000507819523372866,-0.00130635779152333
"3252",-0.00670658616938202,-0.00421952914915569,0.0038779350215703,-0.0051727962225927,0.0209675325407865,0.00891817369642656,0.00609876240846119,-0.0019759370331307,0.00957985388677685,0.000654066522213448
"3253",0.0061702553475107,0.00958965935737455,0.0112529707975328,0.00756330603873012,-0.00998535881126827,-0.00383934588363632,0.00389697467081307,0.00222725231174592,-0.00136584716148491,0.0156862734681336
"3254",0.00179803227216468,-0.00176710696361793,-0.00398610609393146,0.00445691502323831,-0.00486408007566419,-0.00233031240946091,0.000862637697785607,0.000987548869418653,0.000575885409960897,0.00193043642338497
"3255",0.00913410709482765,0.00885142570053654,0.0115057694300502,0.00583836257087689,-0.00553447784262417,-0.00305449840201233,0.00172377718564931,0.00666022259127996,-0.00992809352517998,0.00642265108196249
"3256",-0.00314427453402788,-0.00438683764496306,-0.00560502758531856,-0.00394708469700766,0.00216817640013689,0.000810924103102906,0.00204339791576502,-0.000980261927361004,-0.00029060457384833,-0.00127634574400448
"3257",-0.00111512918704404,0.000440569178826955,-0.000497333434168246,0.00349646593713482,0.0000723740013319762,-0.00117033812329204,-0.00601047243854536,-0.00171687972179868,0.00283470703830924,0.00447288663458867
"3258",0.00283876293987761,0.0048448502773053,0.00215617256771994,0.0146341584549416,0.00786102763571184,0.00414657727766876,-0.00971828551748266,-0.00196563429450769,0.00688553303699702,-0.00445296900902392
"3259",0.00861905937815921,0.00832775356032411,0.00248267031145954,0.0173992551920621,-0.0164581191081163,-0.00790017663595377,-0.0130846422156485,-0.00467746464010688,-0.00352724594770004,0.00894570834782171
"3260",0.000599135317791655,0.00912848508098341,0.0026415535094968,-0.000450009046657818,0.0115679287976458,0.00588184903713351,0.000994343484978399,-0.0029680740933401,0.00447887041358164,0.00506645466891054
"3261",0.00686997784289911,0.0133553272715339,0.00459903204203194,0.00848460157239006,-0.00899041888592844,-0.00467775106171164,0.00642051375819275,0.00620199952358136,-0.0000719884917945723,0.00693133829067927
"3262",0.00021922199845803,-0.0070603627388407,-0.00215629631222214,0.00911985583204378,-0.00137868692246368,0.0000903205823488129,-0.00852825710827998,-0.0066569372801798,-0.000215750873923115,0.0043804543080963
"3263",0.0000625639267366473,-0.00107732450898435,-0.0039893627310138,0.00542253031209938,-0.0082124033892419,-0.00271151347020515,0.0129581084205801,-0.000992723425900066,0.000072002016833439,0.000623031858375089
"3264",0.00409900532174268,0.000215684078000766,-0.00100127204494405,0.000449434712705754,0.001599890729723,0.000780548829576233,0.00827088318189695,0.0084471599886824,0.00258956257834675,0.00435869731147753
"3265",0.00438415809173365,0.00345044303798581,-0.000668262617268822,0.0020215590663426,0.00131887719648005,0,0.00623427239037144,0.000985467132060824,0.00100444106025099,-0.00123988358548832
"3266",0.00152776756569195,0.0023641418488618,-0.000835836116578115,0.00134491114121515,-0.00146343778358238,-0.000906660828253081,-0.00565211463144832,-0.000157303878370874,0.00308194515246707,0.000252270433905188
"3267",0.0000311640518946277,0,-0.00401546097139127,-0.00223859897063661,0.00285808385498654,0.00172432436072434,0.00273281718006513,0.00262193709928171,0.00943199019861352,0.00441361916771754
"3268",0.00532318504189888,0.00385933424576312,0.0026877326067094,0.007179753087174,0.00241175853897269,0.00144968505638632,0.00534179961539172,0.00679919860374878,0.00785730139853325,0.00753289391086009
"3269",-0.000247782697829324,0.00384449704665313,-0.00184273590032824,0.00400983856082804,0.00109358742138022,0.00144765967447524,0.0027108882225082,0.0064933767775861,-0.000351193975586694,0.0018692213002629
"3270",-0.00551315262736363,-0.00680849344448553,-0.0088957179571485,-0.00665628309712052,-0.00364097181867962,-0.000632489778020884,0.000757015280203666,-0.00206447196973514,0.00210779874787059,-0.00186573383084565
"3271",0.00242925450533171,0.0059982791456783,0.00321768664351008,0.00223350763999197,-0.00979422262851926,-0.00361591683265183,0.00583531450190677,0.00310320730784053,0.00189293269673496,-0.0062304676779108
"3272",0.00935184405578715,0.00787915157836161,0.0104659135570777,0.0202808251531668,0.0112933373108448,0.00462701435214163,-0.0110657739472768,0.00206242247327992,0.00734781696351927,0.00125391849529799
"3273",-0.00757211560282867,-0.0107755068864567,-0.0110257753415084,-0.0185669723319049,0.0154004259862184,0.00668314696807015,0.00716990463969425,-0.00205817764145821,0.0132685240695074,0.0118973074514714
"3274",0.00381503979291264,0.00363101916410558,0.0035472874833693,-0.00244833554007728,-0.00567846850130227,-0.00107679502548697,0.000863031856573215,0.00232027829556136,0.0104894967058171,0.00185649752475237
"3275",-0.00281184001572976,-0.00574600153729676,0.00168319177431009,-0.000669350219466014,-0.00491597032789759,-0.00143685373740565,-0.0101305205418367,-0.00360093716501375,0.00393515166520908,-0.000617726953815456
"3276",0.00532965494710136,0.00192639568344166,0.000168065246451743,0.00580489050953625,-0.00661075611874629,-0.00233844363609914,0.00239519495736529,-0.00722755651930396,-0.00750152052779929,-0.0148331273176762
"3277",0.00678051155553705,0.0029908103632359,0.00705643216125584,0.00665921603219544,0.00351032477167035,0.000721361130259668,0.000543197507445914,-0.00078017813394593,-0.00565165459858608,-0.00439146800501888
"3278",-0.00287767467021516,-0.00489885064817175,-0.00700698782699993,0.00529231064326297,0.00889062989417355,0.00216188602558431,0.00868425042351628,0.000520515939787414,0.00602619328922938,0
"3279",0.00687731098311506,0.00449485777111458,0.00571242513457548,0.0155735024638237,-0.00303366423556062,-0.00116842313268828,0.0106543217444832,0.00546165144821487,-0.00741948791996483,-0.00756143667296783
"3280",-0.00152456126425338,0.000639258518361441,0.000334080595595587,-0.00561548542336943,0.00514400447835039,0.0019799300163712,-0.00383347987053484,-0.000776035686098964,-0.000891544326973026,0.00444444444444447
"3281",0.00225981229406313,-0.000638850127975266,-0.00367401412599566,-0.00781933701297721,0.00663172822352509,0.00251475326698136,0.00887226004640462,0.00336521119964783,0.00583424386252673,-0.0050568900126422
"3282",0.00831838222603221,0.00554013183047131,0.000670485914274987,0.00634851785087265,-0.00315096957538608,-0.00206066117170312,0.00741689923623601,0.0064499262945148,-0.00156950328228833,-0.00127064803049548
"3283",0.0031126961432304,0.00487393625989374,0.000670053613780919,0.0056558850142765,-0.00854796660117796,-0.000807967705902413,0.00115695123230308,0.00410150373710394,0.00184542412474098,0.00318066157760799
"3284",-0.00195824588417848,-0.008013496424086,-0.00535667015753771,-0.0253082535692041,0.0105053323646671,0.0039532291807145,0.010190093896105,-0.00663774191197808,0.00109157455189557,-0.00570703868103994
"3285",0.000120672834161839,0.000637763661286872,0.00454393659567898,0.00821126653488236,0.00351356479117104,0.000179107615461582,-0.00571964682651882,0.00411215051067537,0.000340656932647843,-0.0133928571428571
"3286",0.00114689615444474,-0.00403650878987383,0.00117268864678199,-0.0103456294581246,0.00700174264444198,0.00250537527360484,0.00596177921148855,0.00204764183152695,0.00224812327635981,-0.0084033613445379
"3287",-0.00889309053173137,-0.00234640426539845,-0.00384870338005205,-0.0080071009283702,0.00808880997093775,0.00357008818146487,-0.00228744926807634,0.00229894228327554,0.00584557523944995,-0.0149934810951761
"3288",-0.0160293879559114,-0.0205260126986779,-0.0179741183180622,-0.0345290635558105,0.0155544073544636,0.00675915045972286,-0.00479360723293598,-0.0127422635106216,0.00682530765847567,-0.0185307743216413
"3289",0.0104791248533731,0.00873167914856721,0.00889499364190804,0.00836029120447934,-0.00783114055095957,-0.00335677838000237,0.00429309501713626,0.00129067774754521,-0.00892678002125047,0.00472016183411994
"3290",-0.000826043077930771,0.00129843770774341,-0.00322136821414076,0.00483661928695156,0.00977909096419127,0.00478615336971866,-0.00312787916638446,0.00567150276215589,0.00541787199193089,-0.00469798657718123
"3291",0.00324542542171669,-0.00129675395351248,-0.00136085049782564,-0.0148980875188839,0.000138510245854873,0.000970537181955278,0.00125515279901611,-0.000256269854291502,0.0000673177928653956,-0.00876601483479433
"3292",-0.0181579282385191,-0.0157974380674126,-0.0163515457464531,-0.0202419465505873,0.00912973380950666,0.00502326189816449,-0.0121174282291575,-0.00410255509830115,0.0057924226726449,-0.00816326530612244
"3293",0.00742860975456416,0.000879564140558786,0.00761901164058587,0.0111612180961322,-0.000810150055933323,-0.0008516118192059,0.00306650989170909,-0.00102993664695727,-0.00649568731673889,-0.0185185185185185
"3294",0.0152411337699194,0.0158172555271905,0.01512294158899,0.025833787517118,-0.0134668814004519,-0.00580026450262194,0.0102256304387891,0.0048970176752936,-0.0130089511120994,0.00139762403913335
"3295",0.0115480788669458,0.0114619142142474,0.00897231702770407,0.0057234102491881,-0.0109346544753313,-0.00433121194161323,0.00020858827874215,0.00051282892436344,0.00122931099231849,0.0153524075366365
"3296",0.00336483736673454,0.00171039020727148,0.00755039526441625,0.000910486163524959,0.00450652263346996,0.000710209616109347,0.00375596571140902,-0.000512566065659414,0.0053883977533018,0.00412371134020617
"3297",-0.00532968105364606,-0.0087512560463181,-0.00965854307418046,-0.0138730461421211,0.0124781188464527,0.0047906716027506,-0.000415849981605376,-0.00461664699596231,0.00264585492452607,-0.00547570157426425
"3298",0.00746539614223063,0.00258401394480279,-0.00117709476595496,0.00553501241271737,0.00276943215010128,0.00194241842979892,0.0100863299096539,0.00566868613223792,0.00257124986804746,-0.00894700619408118
"3299",0.00173299510010061,0.00601367272510611,0.00505051038477689,0.0130733985207427,-0.00504013085813149,-0.00237932479716951,0.00813257347395657,0.00358688754167891,-0.00344195185856722,0.0034722222222221
"3300",0.00644282192660373,0.00576440322925542,-0.00485766835444512,0.0135839826710751,-0.00506609135163882,-0.00256174933810649,0.00796482119314956,0.000510682356676728,-0.000812752246708404,0.013840830449827
"3301",-0.00106699100346452,-0.00785399861214608,-0.00875275733086789,-0.0131785349111432,0.00383619208365515,0.00088571506960311,0.00678755194453129,0.000255223964669593,0.00569345289314205,0.000682593856655256
"3302",0.0016021507004127,0.000855787658175622,-0.00747145325008181,0.000452759021563942,0.00437732484399977,0.00247746100788326,0.00905616004558607,0.00867343342949622,0.00417842687092507,-0.000682128240109159
"3303",-0.00257705704258804,-0.00448909259205321,-0.0148845560352959,-0.00656118412657902,0.00684891276378363,0.00158873661172398,-0.000697903515503917,-0.0035406226365815,0.0128188187919462,0.00750853242320826
"3304",0.00478115848824401,0.00579767003434917,-0.00173675697544018,0.00728764697794615,-0.0000687234249293622,-0.000176320411576114,-0.0125736984590221,-0.00304581523019831,0.00583121712726231,0.00948509485094862
"3305",-0.00410806239924344,-0.00597772464544755,-0.00643702394936052,-0.015600208138483,0.00783344245690532,0.0029086031740031,0.0108135001576675,-0.00381877636813255,0.00408466320964895,-0.00402684563758393
"3306",-0.0102983128434405,-0.00279211162313076,-0.0084048172260508,-0.00574183682717067,0.00934076885989921,0.00404252928778015,0.00189976625999844,-0.0020445021867882,0.0150252144865768,-0.00404312668463613
"3307",-0.0331654841572129,-0.0432910056289861,-0.0337276689080698,-0.037422120924021,0.0149284025253182,0.00778980354538339,-0.0133719020933517,-0.0197183324066023,0.00898512622466319,-0.0189445196211095
"3308",-0.0303021541737136,-0.0229625929431726,-0.00164475335735925,-0.00791931751893882,0.00532432059349963,0.00277920035940671,-0.0268029471572216,-0.0107104156142139,-0.0178742588986933,-0.0186206896551724
"3309",-0.00367809893143067,0.000921553809988707,0.00494233351506534,0.00798253373821733,-0.00529612234025767,-0.000519558026391143,-0.0104967451463084,-0.0105624948312235,0.00437050219757662,-0.00983836964160234
"3310",-0.0449116854613356,-0.0303867507086837,-0.0342440848056547,-0.0239980900206995,0.0108485642562677,0.00485267082957774,-0.0524103895322263,-0.0240192967046704,0.000194836655226238,-0.0170333569907736
"3311",-0.00420163344118829,-0.00807208989720432,-0.00113167255195179,-0.00368815636707587,0.0225834544298946,0.0112108346295077,-0.031257029296289,-0.0213287903680033,-0.0364934740259739,-0.0173285198555957
"3312",0.0433064257416271,0.0179512180975343,0.012651142624619,0.0217176519164763,-0.0073571912081476,-0.000683148761897345,0.048169318376073,0.00558810451230629,0.00552629715843445,0.0227773695811904
"3313",-0.0286322964268988,-0.00893489292641636,-0.0128660557251218,-0.00676335529423111,0.0155255875767066,0.0116200553229637,0.000109261450937925,0.0133370084178119,0.0314343303907707,0.00215517241379315
"3314",0.0420329259550256,0.0360616346656353,0.0217227742669746,0.0177528930520168,-0.0106186356008368,-0.00219599675309301,0.0382012244533574,0.0235811182574088,0.00175453246965063,0.000716845878136363
"3315",-0.0332416353354782,-0.0316005984418652,-0.0181179385232649,-0.0210273908471711,0.0248916268941317,0.00888785378084833,-0.0217620450391843,-0.003750426128449,0.0216009400207333,-0.0107449856733525
"3316",-0.0165310689540706,-0.015133562716705,-0.00960278247085289,-0.0205028464407714,0.0520439767081853,0.0101519213701489,-0.0169800680998408,-0.0188221709390026,0.000380963858627181,-0.0325850832729907
"3317",-0.0780945347457551,-0.0871548986612232,-0.0509505688500164,-0.0682780508424983,0.0271031794684842,0.00896993973442517,-0.0741227561632529,-0.0570019851747433,0.00165023798825326,-0.0778443113772455
"3318",0.0517449123039622,0.0360336123254741,0.0298477995090447,0.0508158210399736,-0.0512579593830528,-0.0183568847646953,0.038611429945997,0.00610286167445473,-0.0211013373183111,0.0316558441558441
"3319",-0.0487483516908587,-0.0558517127924183,-0.0338455487657232,-0.046576875817241,-0.0367978705355492,-0.00997909846671186,-0.058208287207507,-0.0283073450178859,-0.00356035094666884,-0.0180959874114871
"3320",-0.0956772442428522,-0.113471321790685,-0.098047109369466,-0.100106782456036,0.00619686503200012,0.000508294964395306,-0.0974167629323441,-0.103448270592329,-0.039888262711738,-0.0400641025641025
"3321",0.0854862023186675,0.0606612444536092,0.0328124991882823,0.0720854973569889,-0.022603113449759,-0.00651875906661226,0.0853285263816004,-0.0135941920931343,-0.0305162339374359,0.0108514190317195
"3322",-0.109423646457338,-0.113239970988953,-0.0659174392301433,-0.124792503442331,0.0647655522431234,0.0264166453420316,-0.168699956403489,-0.0988234920045739,-0.011446119566207,-0.060280759702725
"3323",0.0539920388008523,0.0451467391865614,0.0490513725951562,0.0689219232106981,-0.066683036412123,-0.0250727050033148,0.0469907171376105,-0.0193957337079046,0.013555485834196,-0.0158172231985941
"3324",-0.0506329488316828,-0.0688059631979527,-0.0211733393062021,-0.0863650036482236,-0.0564126370322249,-0.0138805683128341,-0.0984000068590882,-0.0928109729441079,-0.0199219910827807,-0.0330357142857142
"3325",0.00212495995971218,0.0218687765267744,0.0139702730661881,0.00776951055149566,0.0272255818697908,0.00328154096918376,0.000471032755124501,-0.0612159433256795,-0.0189055014692003,0.0212373037857803
"3326",-0.043094127850326,-0.0126458857656078,0.00244437651511475,0.00738842855908461,0.0751956363200998,0.0254777506754045,-0.0437922112360217,0.0236713647440396,0.0149957121484352,-0.0108499095840869
"3327",-0.025568229035413,-0.00821015664447389,-0.0104189439520959,-0.0239158409604547,0.0412091614661867,0.011834792448268,-0.0505580865176194,0.00334731273147448,0.0441795871516695,0.0118829981718465
"3328",0.0906032779960004,0.0894039533811828,0.0694445036328,0.0751388918214073,-0.0186144424737293,-0.0068021989403354,0.0800484551109599,0.0930640970784973,0.0485303544388853,0.0216802168021681
"3329",0.0149701928235477,0.0407294397318521,0.0188520075776331,0.0352476173013849,-0.00227114312332588,0.000584592055269395,0.0549026180283649,0.0650602512143974,-0.0136896419956835,0.0167992926613616
"3330",0.0583897580537081,0.0487733643902877,0.0328948014432142,0.0378632715921607,0.00492188676755623,0.00242063471223153,0.0741536340838187,0.0282806118894561,0.012822220499229,-0.00347826086956515
"3331",-0.02978565678878,-0.0345308092337697,-0.00119429294900686,-0.0568440936789796,0.0266928480015645,0.00741129679268915,0.00128361432832258,-0.0352036366302383,-0.00646048660726684,-0.00349040139616064
"3332",0.0324757391536492,0.0187482439645701,0.0121562211409505,0.0164919182175003,-0.00822907589038402,0.00231436573260901,0.0199430959073672,0.00836199565726536,0.00440064367816095,-0.00262697022767067
"3333",-0.014905338203151,0.000283187261510998,-0.0275645048702315,0.0067846830326328,-0.00811692421463206,0.00181426527719197,-0.0283519315480202,0.00904629620280839,-0.0318466849574507,-0.0122914837576822
"3334",-0.0450048893438236,-0.0467024793622237,-0.0475803782906949,-0.0427776690019332,0.0140106824257031,0.00407129924597238,-0.0659767136077433,-0.0362346586816086,0.00945622405694913,-0.0284444444444445
"3335",0.0230754164745575,0.0190023559480119,0.0127549644120442,0.0336700222543904,0.00634599835507288,0.00016403534216014,0.00430911891221686,-0.0104650852944225,0.0163934228784226,0.019213174748399
"3336",-0.014454203616645,-0.0203963939590336,-0.0224600386189324,-0.0189516763023175,0.00237932504993044,0.000738831404663909,-0.0156298788909269,-0.0336857722805298,0.00493745904953746,0.0251346499102334
"3337",0.0671661852708443,0.0475908451064415,0.0590508819167488,0.0546332215093448,-0.0026113447973658,-0.00451053609697427,0.0750311641473511,0.0381029516962397,0.0277105218883926,0.00525394045534155
"3338",0.00101949519586308,0.00454293401315931,0.0107461236419419,0.0051517069219118,-0.0104724565939451,-0.00444830981300703,0.00970173943394648,0.0394376513755572,-0.00535448733571875,0.00696864111498252
"3339",0.0335684049000033,0.0146975627787778,-0.00240725273821429,0.0102505478571475,-0.00727594746066063,-0.00124142472612188,0.0715616620871093,0.0202855150895977,-0.00890796630579194,-0.00259515570934266
"3340",0.0152172750358999,0.02395535252479,0.0130706705692862,-0.0036641079871883,0.00181700546660801,0.00215427612053753,0.0556744959554432,0.0261414303111067,0.0261235574312406,0.0026019080659152
"3341",-0.00913008716805042,-0.0141457223873751,-0.0041683893940716,0.00141451693496375,-0.00912969164658706,-0.0021496451912344,-0.040694789627386,-0.00717616525115194,0.0171403488923014,0.0173010380622838
"3342",0.0294928734580193,0.0187636521564496,0.0183376939379931,0.0228813077641175,-0.000244176560704745,0.0013255947800892,0.0264306214200554,0.00542098010660719,0.00786809347950945,-0.00850340136054417
"3343",-0.0212480717679999,-0.0392740533355447,-0.00998239870540929,-0.0256834974030193,0.0264891608634084,0.00893614225427419,-0.0378523208621818,-0.0287562888330475,-0.00510196112437744,-0.0205831903945112
"3344",0.00482424045424024,0.00281920658165657,-0.00850139186469856,0.00538546035734333,0.0113571622430837,0.00106599457325074,-0.0112405497883554,-0.0074019146513068,-0.000864992244733132,-0.00262697022767067
"3345",0.0270153491771443,0.0334552359857732,0.0133599295051732,0.0222723290695688,-0.0134049300173702,-0.00262136063781415,0.0297738002027301,0.0294556039319709,-0.0194174748876239,0.00438981562774354
"3346",-0.017617918356675,-0.0136018119398276,-0.0153482967970563,-0.0126861982538108,0.00804481854933847,0.00262825022951207,-0.0362726429116983,-0.0130387516830515,0.00712612694782822,-0.0166083916083916
"3347",-0.0303632409252813,-0.0206838898200327,-0.0093925380970391,-0.0276533775518809,0.0125917175817625,0.00278532922441932,-0.0182736018241177,-0.0264219386860173,-0.00682527251393739,-0.0471111111111111
"3348",0.0221945517829849,0.0152069289882333,0.017349220352503,0.0272908074199041,-0.0102167560753946,-0.00310442156172652,0.0159744283097718,0.00980013182525785,0.0196708592165005,0.0139925373134326
"3349",-0.0000717539684833568,-0.00776698150173061,0.00138803881588667,-0.00363519088247444,0.00530857944710439,0.000655759264749367,-0.00916054360385465,0.00373271221196769,0.00995486328955342,-0.00275988960441576
"3350",0.0139388175704263,0.012300833365315,0.00772289741842513,-0.00140337209165364,0.00234693227686233,0.000245455793644211,0.0041396494715995,-0.000371833849167391,-0.00428552110409031,-0.0129151291512916
"3351",0.0144184624209178,0.014360697385033,0.0137551591142424,0.0202360155888257,-0.0186136401213581,-0.00532169154765905,0.0316064915865553,0.0171131065150638,-0.00664043904722345,-0.0186915887850466
"3352",-0.00459855883267413,0.0070787214817376,0.0145376964703137,0.00192831776432723,0.0115111727692458,0.00436250066460087,0.00905812501039449,0.00658377728160797,-0.00445656108512704,0.000952380952381038
"3353",0.0261785484847687,0.0267638511312289,0.0175772628270587,0.0291449275755107,-0.00518903254886083,-0.000491653405560233,0.0153136210991232,0.0243458804204391,0.00553344952831258,0.0180780209324451
"3354",-0.00931062168673058,-0.0184307598014206,-0.0281637384778045,-0.021106051525421,-0.0116768155899956,-0.00237784326105162,-0.0111818769721779,-0.00638525989898464,-0.0181165712759925,0.0186915887850467
"3355",-0.026473529743954,-0.0206544840774022,-0.0175810573075463,-0.0360262559189392,0.0085633992610703,0.00138221183293585,-0.0339251099502293,-0.0199928483209154,0.00617125932925822,-0.0128440366972478
"3356",0.00275833719416552,-0.00109546532665772,-0.00491645266148966,0.0107589247284108,-0.00470383757720072,0.000164462416771149,-0.00299438542493535,-0.00546446445131643,0.00350480037241718,0.0120817843866172
"3357",0.00923924808653598,-0.00219366895985551,0.00968382784631361,0.00560225413218629,-0.00640101334927856,-0.000739467452362086,0.00477816767120709,0.00366294285011515,0.00424103790048735,0.0257116620752984
"3358",-0.00677866164862895,-0.00741963630183418,-0.00763363163184849,-0.00306405706733404,-0.0161358430993236,-0.00369940343951958,-0.016576189940629,-0.0113137855469899,-0.0128555890484265,-0.0196956132497762
"3359",0.0120667804285479,0.0166113777638426,0.0149901654656659,0.00810285801088462,0.0167062810302516,0.00610610549619151,0.0132633475877055,0.0184569515255051,0.0153507520984728,0.00639269406392695
"3360",0.0165462030750507,0.0166121446208018,0.0171007173751914,0.021064276852909,-0.013000899757725,-0.00328055760915058,0.0238613415257125,0.0224718918619804,-0.00601029187688384,0.0208711433756805
"3361",0.000205127339911071,-0.00482184181478107,0.00955290730397929,-0.006514717281914,-0.007805875259836,-0.00279766755383182,-0.0141162440767205,0.00248151455427492,-0.00623363678136934,-0.0133333333333334
"3362",-0.0199315157701656,-0.0123823177141621,-0.0130583565157129,-0.00382524569981924,0.0102642994891142,0.00330058903999819,-0.0459273411170292,-0.0275814238776146,0.00388906666527511,-0.00810810810810814
"3363",-0.0176859348775098,-0.0136276528142779,0.00479389508967598,-0.00191985570952902,0.00699631667587886,0.00205615012795102,-0.0236442875409159,-0.0152727923759035,0.00962265100823889,-0.0099909173478655
"3364",0.011967419914134,-0.00828952510127301,-0.0148855046520197,0.00384720899184843,0.00978742358809725,0.0015593757813579,0.00464037613741453,-0.00443126395712379,0.00885006177930348,0.0174311926605504
"3365",0.00459698385030394,0.00167171199142113,0.0017435278612099,-0.0136873302113096,-0.00257271910292522,-0.000655695863170491,-0.00461894250682571,-0.00964390060318909,0.00564381343610254,0.00991884580703339
"3366",0.0304595666041756,0.0445062614152016,0.0249468417981387,0.0391339059951523,-0.02195428109377,-0.00614993635900374,0.0582946873223136,0.033333321889516,-0.00756414965502994,0.0285714285714287
"3367",-0.0102711891870366,-0.0143808831070626,-0.0116981268387597,-0.00801267797322114,0.00374118593109651,0.00280528495907939,-0.0112359308712536,-0.00144982090979595,0.00965021194111237,-0.00260416666666663
"3368",0.0169880592511369,0.0224265087330278,0.0150819758905292,0.0131933431690099,0.00299390068006855,0.000246670327197718,0.00970060166341979,0.00725959274279542,0.0023742786550065,0.0174064403829417
"3369",-0.00690391241473809,-0.00845666486189389,-0.0107202752048039,-0.011427058373339,0.00249776291805337,0.000658243204793685,-0.0013724362947134,-0.0100901205235654,-0.014576338217176,-0.0042771599657826
"3370",0.00189911727406167,-0.00266525366460491,0.00133077561348682,-0.0206989411435453,0.00601614847385812,0.00189058410898291,0.0136062984964016,-0.00327632861658333,0.00591683821263467,-0.00773195876288657
"3371",0.012320455604274,0.0253874787444441,0.0339851812722056,0.0219599478036063,-0.0134097977825437,-0.00262558227837129,0.0364746727305048,0.0365229995509746,-0.0142148636756079,0.0103896103896104
"3372",0.0148790539888781,0.0138129533654103,0.0128535472905713,0.00322312738288866,-0.00183684946453921,0.000822714409023817,0.0192307471612778,0.00845670620548811,0.00180243645846501,-0.012853470437018
"3373",-0.00184499958864637,0.00925435979006495,0.0130529400635941,-0.00696109714413318,-0.00368035417484236,-0.000904174937475299,0.00410721584351048,-0.0027952514852676,0.00335034137890799,0.00520833333333348
"3374",0.00445597019512034,0.000509457183774931,-0.00841092697984491,0.0172552725783459,0.00714157552262451,0.003208594230804,-0.0103540560578326,0.00875970429676975,0.00735841573486007,0.0172711571675301
"3375",0.00404165392613964,0.0224033257097773,0.0151597501810032,0.0230585436619108,-0.0067328621720536,-0.000394148442928399,0.0231207302634346,0.019451150029032,0.00460376883914382,0.00594227504244493
"3376",0.00828007398306752,0.0114541585033494,0.00444440135024293,0.0238342236541351,-0.00363568013910265,-0.00164240039709185,0.00896344995513032,0.0252129514573673,-0.00647682985514275,0.0109704641350212
"3377",0.0133083942407244,0.0295420660014845,0.00690269497532525,0.0232794034716983,-0.0132968646196531,-0.0059225518554481,0.0300300170751049,0.0312396095852701,-0.0184501838210265,0
"3378",-0.0026267616300476,-0.00310850464199064,-0.0112497772418638,-0.0140949587704999,-0.0144793647293332,-0.0039718084760022,-0.00850333377805279,-0.00902352005641893,0.0105262715341001,0.00834724540901499
"3379",0.0256294639269152,0.0191892656951858,0.0144000193995864,0.0263355767654689,-0.00712315043051404,-0.00498462510068265,0.0363880293353076,0.0198373600063886,-0.02027532254635,0.0198675496688743
"3380",0.0120875439359664,0.0115320150753384,0.0147213582776899,0.00610947167774101,0.00384358994515233,0.00108551541113178,0.0263623933244534,0.0191325954796409,0.0108221381818283,-0.00649350649350655
"3381",-0.00745668151774781,-0.0155885234072978,-0.00518142258028087,-0.00680106531000779,0.0113583778945909,0.00358626106670279,-0.0161252841610054,-0.0134542038069074,0.00964183565212973,0.00326797385620914
"3382",-0.00557997223741902,-0.00354533253245415,-0.000520774198199847,0.00733662561794324,0.0148273256734988,0.0074794478364022,-0.0255209745103122,-0.007294757617751,0.014324767900433,0.00651465798045603
"3383",-0.0576489166702419,-0.0600094210254433,-0.0420357413269354,-0.0521970203829051,0.0189009267750695,0.00354698309919432,-0.0631906206152847,-0.0578274572836955,-0.0072140854038113,-0.0323624595469254
"3384",0.0119756321599045,0.0181678849337092,0.0179510392575122,0.0212602762118725,-0.00964123144022422,-0.00221936642260723,0.0357782149064969,0.0267887890148186,0.00141631874756021,0.00418060200668879
"3385",0.00933562742433436,0.00963484717817509,-0.0109160742471491,-0.00908183101356075,0.00055445973703705,-0.000823795675292116,0.0115035887298527,-0.00825630592771898,-0.00178325549696379,0.00915903413821817
"3386",0.0192477277485787,0.0119283280385221,0.0192412739727763,0.00636464387278179,-0.0153334672389865,-0.00206107118113641,0.0197140936469109,0.0116550220907274,-0.000492835575767514,0.00825082508250841
"3387",-0.00415395001656094,0.00319255550010489,0.00445237772557805,0.00961298798860222,0.00412767416072901,0.00156968944364255,-0.013533167557409,0.00592489935526097,0.00191061941448378,-0.0049099836333879
"3388",0.000385058377969427,-0.00758870775860954,-0.00177312441225086,0.000501118726354832,0.0105879831696425,0.00222711412609655,-0.0106564668349824,-0.00589000168805687,-0.00196846090020264,0.00575657894736836
"3389",-0.0057148570425456,-0.00370012522609997,-0.00479574177844944,-0.000250471820186893,0.000801059526321257,0.000329229865733138,-0.0126284299153128,-0.01547066925223,0.0110330001530756,0.00817661488143906
"3390",0.00641517217094179,0.0143600662384726,0.00678214537879995,0.0122745236306188,0.000123179467563794,-0.000905046939671528,-0.0018809201310892,0.00752692060578486,0.00646221426850113,0.0105433901054339
"3391",0.00460366655181232,0.00585788303787171,0.00265911728461288,0.00965106995117404,-0.00683451410763813,-0.000329427925807924,-0.00301506961958398,-0.00435514477014409,0.00841965009194134,-0.00481540930979141
"3392",-0.0255086744417172,-0.0266925372598709,-0.0208628035094219,-0.0132352605052479,0.0107252827711779,0.00189483271509183,-0.0286038157624885,-0.0211978679724223,-0.00348391406736948,-0.025
"3393",0.0107204962094321,0.0157068830781257,0.0113759038541403,0.00422259226138988,0.00288306955052064,0.000164361593787632,0.0123232823865629,0.00446892674177124,-0.00060271852692162,0.00909842845326714
"3394",-0.0237513840143926,-0.017918632329166,-0.00964107291646166,-0.0121197873986137,0.0107033092598938,0.00271291693456055,-0.01986171507072,-0.0102669588847596,0.00446314829077532,-0.012295081967213
"3395",0.0146974679067127,0.0119970768093913,0.000180207403029486,0.00450675713808302,-0.00314690768963255,0.000983834170845022,0.0186953737665208,0.00242046883942448,0.000540482789620489,0.0165975103734439
"3396",0.0128095224492002,-0.00222273210838231,-0.0100937048991532,-0.00324018467637377,-0.00485646023668085,-0.00180188202768572,0.0114219927136583,-0.00586407271135569,0.00444091686848336,0.00489795918367353
"3397",0.0070048546154069,0.00816823988803539,-0.00200291924977958,0.011252754144756,-0.00194191372197305,-0.00156051642742649,0.0224590776126579,0.0156141323850161,-0.00448108993490737,0.00812347684809089
"3398",0.00550689525659886,0.00932978087425207,0.00656809568525318,0.0227497784450741,0.00104017449267535,0.00123382394759597,-0.00310255568749196,0.0143492235632483,0.00216061103590848,0.00402900886381952
"3399",0.0154374048655805,0.0184868852878821,0.0128693782473652,0.04303670300978,-0.00409555436313036,-0.00147883349645472,0.000124440525363312,0.00707298211016538,0.00598874131006677,0.00802568218298561
"3400",-0.0103138172182856,-0.0157630259524023,-0.00894772743392935,-0.0166898356743294,0.0140561369266137,0.00320881029486753,-0.0190439684295641,-0.0170568374208426,0.00631025732373525,0.000796178343948961
"3401",0.00764855548698606,0.0111622853159155,-0.000722309247590536,0.0259312101475135,-0.00399516379173703,-0.00155815150390404,-0.00101509759177998,0.00510387204307716,0.00621156556720881,0.0127287191726333
"3402",-0.00569297081568332,-0.013918839964588,-0.00487891663208373,0,0.0159223027983428,0.00320348062766773,-0.00558880637095649,-0.0135410306842894,-0.00270439773542008,-0.0117831893165751
"3403",0.0102106510138127,0.0109515989679205,0.0130742445956868,-0.00643380332254151,-0.00502496455950718,-0.0019650187898802,0.00281015363748827,0.0061770874471303,-0.00259389840848034,0.00635930047694755
"3404",-0.00865898593093406,-0.00481463843321106,-0.00519803705289312,-0.00670678688260207,0.00330681838300784,0.00106643037630905,-0.0123551329810793,-0.00920873072510819,0.00124116081043613,-0.0102685624012638
"3405",0.0129590396870023,0.0164489616254091,0.00792791504741186,0.00139692516972678,0.00143805521482143,-0.0000818703894057693,0.00760891038304568,0.0103270410843739,0.00466356569056314,0.00478850758180371
"3406",0.00918720566984388,0.0128510380881499,0.0126922337458115,0.00302255868954138,-0.00466717133998962,-0.000327870476809045,0.0103674642702687,0.00306642783482847,0.000881332617882036,0.0119142176330422
"3407",-0.00329338927829315,-0.00469924994452819,-0.0102383929563679,-0.0141399606352092,0.00474934264589466,0.000737802342174465,-0.0108944210732403,-0.012228282939188,-0.00945168508751182,-0.00784929356357922
"3408",0.00289900660510445,0.00661000726451766,0.00160515586470078,0.00564309512097294,-0.00209426681677538,-0.00024571166551679,0.012551097844866,0.00412662438045808,0.0082380076628461,0.00158227848101267
"3409",0.00808156825280193,0.00633208976020105,0.000712277195510147,0.0128593847088865,0.00245832346116326,0.00065551831330124,-0.0118895829369681,0.00102727813342107,0.00482016825829334,-0.000789889415481859
"3410",0.00212760332959983,0.00302959330158026,0.000533760675325068,0.00923375202207621,0.000598242722725573,0.00106463251257316,0.00256016533822301,0.00547384999707834,0.0120510002100036,0.0142292490118576
"3411",0.00569205491444502,0.00302037236950059,-0.00266755817373754,-0.00434595694696915,0.00298867320049734,0.000327319314612717,0.0153217140233595,0.00544408441028921,0.0152023410404625,0.00623538581449723
"3412",-0.0119317699176867,-0.00833900223066475,-0.00338805793670549,-0.00804039552719715,0.0116812074245485,0.000981275328810094,-0.00515596876557156,-0.00913705514434771,0.00882530294296791,-0.00232378001549183
"3413",-0.00644037175137901,-0.00700778145068881,-0.00107353232064267,-0.000926385334135249,-0.000058713962867607,-0.000490189499578797,-0.00758426587422745,-0.00102464368324284,0.00857886928576646,0.00155279503105588
"3414",0.0072924215903718,0.0098800133440422,0.0198817545068977,0.0155308973746962,-0.00371166607802997,-0.00155298698928552,0.0115908070717059,0.00649576722463752,0.0197537720160119,0.00930232558139532
"3415",-0.00634237346982991,-0.00372696617641088,-0.00614678988209716,-0.00821729585848896,0.00691856857840456,0.00237415568390809,0.0178795834531074,-0.000339703083125031,0.00834112952513033,-0.0053763440860215
"3416",0.0122987473510801,0.0114566188788765,0.000530099921910443,0.0161104674450836,-0.00170299045483213,0.00130671203206068,0.0223900003452073,0.0190282259851782,0.00751023129251704,0.00540540540540535
"3417",-0.00356794752528644,-0.0147943291059862,-0.0150123321544426,-0.0126840832527064,0.0065885074743437,0.0013865471640615,-0.00508165663462812,-0.0103367583990788,-0.00740025907739816,-0.0115207373271889
"3418",0.00790221208660902,-0.0213514550800794,-0.0258202853673972,-0.00688226131496184,-0.000642867095253741,0.000244478780596191,-0.00206740950299056,-0.00707550136036739,0.00908793015585352,0.00543900543900544
"3419",0.0069521638024781,0.0191800854218376,0.0204305959507118,0.00692995507670058,-0.00503483134123683,-0.000489026115615188,-0.0130393516374125,0,0.00113253523123413,0.0100463678516229
"3420",0.00386260061287347,0.0028228948101634,0.0111833606485863,0.0133057330227853,0.00953228948675577,0.00342459587053545,0.0125942151090994,0.0115371546064917,0.0212777258202852,0.00535577658760533
"3421",0.00621093723544552,0.00492610080761691,-0.000713529813938241,0.0108672348183372,-0.00874292290949197,-0.00333167336532059,-0.00378006445277335,0.0110701139480471,0.00928324298292615,0.00837138508371371
"3422",0.00668459206482286,0.00210080353101283,-0.000714057223142661,0.00313544315669989,0.00558610247583546,0.00114146345509569,0.000122539875566874,-0.00464498733666063,0.0132740680447117,0.00754716981132075
"3423",0.000717969792883633,-0.00605638750273174,0.000357256832081987,-0.0205403224060086,-0.00666605379106722,-0.00211748924041666,0.013584547164482,-0.00200000363190678,-0.0158853010257635,-0.0134831460674157
"3424",0.00298883748259282,0.00257796251906162,0.00482143304684457,0.00250742191128173,-0.00447382925548689,-0.00106092984716222,0.00241487712008026,0.00334006436572887,-0.00345895921030315,0.00531511009870922
"3425",-0.00825463718686148,0.00467510725625608,0.00817482716730655,-0.00272846513464009,-0.0118850412078473,-0.00343131910120087,-0.014454418252028,-0.000998687000471676,-0.0536944113708465,-0.0158610271903324
"3426",0.013942350140091,0.022335875567705,0.0211528909464751,0.013451851754932,-0.00909578824318347,-0.00295140188896037,0.00965546711676724,0.0103298692791276,-0.00466820045939531,0.0107444359171145
"3427",-0.00180788390741571,-0.00591708460596674,-0.00120833482588034,-0.00292463995868275,-0.0106889029587345,-0.00205560564055796,-0.0113788341795864,-0.0042875678765647,0.0236180673271447,0.00531511009870922
"3428",0.0000297818059293853,-0.0107601052047512,-0.000172885105389375,-0.00180495411884918,-0.00390678648148657,0.000494385042565604,0.000122485623386348,-0.00364366947016281,-0.00430921830241404,0
"3429",0.00317660541753262,0.00786856164824923,0.00414869315549549,0.0126581645386226,0.00251258790603015,0.00164707247860862,0.00783544017457727,0.00698144624406805,0.0216939144946717,0.0166163141993958
"3430",0.00216041523140809,-0.00045922393560649,0.00344295762916635,-0.00111606309734713,0.00715203904748885,0.0017265455897757,-0.00473764479525374,-0.000330137001859798,0.00900800536193036,0.00222882615156017
"3431",-0.00416377190595141,-0.00321616014884829,-0.00531826598374119,-0.0122905012545017,-0.00625157881094751,-0.00131327169225148,-0.0179421503489544,-0.0142007791234133,-0.0315654597776502,-0.00296515937731656
"3432",0.00311362402447113,-0.00276564312393557,-0.00362193036605207,-0.00316745657070705,0.00903939870442305,0.0028764652256017,0.00907285655711165,0.0130652653216625,0.00691393198765544,-0.00148698884758358
"3433",0.00354730219114585,-0.00924428393270871,-0.00276961962482858,0.00499314937346873,0.00599221262637273,0.000737529700233663,0.00147791809446218,0.0056216756353944,-0.00801090463215259,-0.00967982129560674
"3434",0.010133241227593,0.0158619100292168,0.0111091946087025,0.0110660127272986,-0.00162453127022466,-0.00139212055281401,0.00787118346695936,0.00361730975409325,-0.00565840249221783,0.00526315789473664
"3435",0.0034993040256639,0.00229625847229076,-0.00137342436182752,0.0100513889207965,-0.00765375535851476,-0.00237793124087327,0.00244051406928114,-0.00229360959694436,0.00121547513812148,0.0082273747195214
"3436",0.0100255797081819,0.00801833056688506,0.00275062650110192,0.0026536687370784,-0.00382611388819543,-0.0004110370528424,-0.00937312802762746,0.00591127445966766,0.0118088510550225,0.00222551928783377
"3437",0.00218651158521044,-0.0129546234667604,-0.00925773160886156,-0.0083811738077767,-0.0170088980339356,-0.00353587063285155,0.0142541832988798,-0.0111001613587999,-0.0115619327467172,-0.00370096225018501
"3438",0.00645945018783722,0.00736820979544217,0.00536426261288692,0.0131228269773582,-0.000744258663535335,0.00165033792546976,0.00617884882532849,0.0158467759300682,0.0173802356714787,0.00668647845468051
"3439",-0.00362252408184494,-0.00937142324504048,-0.00137690110974764,-0.0221734124888563,0.00664092788786963,0.00107111381214509,-0.0096328179140005,-0.00682479269209402,0.00238626282545851,-0.000738007380073902
"3440",0.00941855675140468,-0.00115359940494186,0.00275766837334324,0.0170632407409088,0.0114377026541443,0.00327772475112953,0.00109417819682567,-0.00163613409122609,0.00119028836021973,0.00147710487444619
"3441",0.0144639807202169,0.0159389143064579,0.0099690090488056,-0.00264896024351624,0.00952044866041524,0.00139547649926564,0.0182171917520215,0.0114716748243153,-0.0131316290764936,-0.0132743362831859
"3442",-0.0344142688239503,-0.023874475997593,-0.0175289211737244,-0.0190349948756297,0.00284118612565498,0.00131170974392236,-0.0124045446781693,-0.0123137183262474,-0.00810423853094511,-0.00896860986547088
"3443",-0.00816480053810109,0.00232935092694975,0.00554304264397731,0.000451255627045954,-0.0189883709453629,-0.00556702235669049,-0.00458936622229011,-0.00492125225186135,0.00276029591895943,-0.00904977375565608
"3444",-0.0273228876179307,-0.0141761765895759,-0.00826873004272743,-0.0173657674001291,0.00614465212522619,0.00214046844052662,-0.0124969872394683,-0.00527529236653279,-0.00192692139356365,-0.0243531202435312
"3445",0.0197473784058546,0.0238095492544381,0.00347405615827245,0.0149185033495722,-0.00268710868384925,-0.000492944834635911,0.00909200560173051,0.0129267549760068,0.00970825786285956,0.00936037441497661
"3446",-0.0173636608959636,-0.0135850251781845,0.000519254804014935,-0.0160561099279276,0.0050826225793339,0.00123286687288116,-0.0133933661907657,-0.0143979205802336,-0.00322314116542255,-0.0100463678516228
"3447",0.000509075696082162,0.0102707413607641,0.0129757966819781,0.00965296998983645,0.00213244159426318,0.00155980173095438,-0.00555343645047857,0,-0.0000548613373668738,0.00702576112412179
"3448",0.0131713037913834,0.00231058357656111,0.00717335708694722,0.0161621030862584,-0.000060831968378916,-0.000901621163760136,0.026805593221801,0.00830017572705133,0.00789258439943952,0.000775193798449703
"3449",0.00505238838467936,0.00691560870099028,0.00457860355758033,0.0105286812983463,-0.00243183932310687,-0.000492191565250266,0.011602490338402,0.0125122590799907,-0.00239274567617997,0.00542215336948115
"3450",-0.00396865640931066,-0.00114464297171923,0.00354491103286558,-0.00133010344579598,-0.00298672126025634,-0.000574554259447857,0.00537647816830256,0.00910578448927057,0.00283458167622652,0.0184899845916795
"3451",-0.00879518780437549,0.00229197863125852,0.00117744049344926,-0.00399555765073989,0.00305664484540125,0.000328464297799869,-0.0187759619404696,0.00515628776022314,-0.00548999290378871,0.0113464447806353
"3452",-0.0115127660144453,-0.00914706509708973,-0.00436828179729654,-0.00780027642787029,-0.00310821258329963,-0.000903044008685461,-0.0215575068008812,-0.0182751044095527,0.00131170742685871,0.0044876589379208
"3453",-0.0111295572353215,-0.0309254077217416,-0.0148498076477788,-0.0092093977355211,0.00507414080334789,0.00180771223055398,-0.0278499701017606,-0.0254027873875655,-0.0200872983638749,-0.0245718540580789
"3454",0.0101843942287585,-0.00261971065479116,0.00308330215764419,-0.00748126865524301,-0.000790644640078275,0,0.0117137601634076,-0.00202839756592288,-0.00484631228060806,-0.00458015267175571
"3455",-0.0231909946794753,-0.0126552295240323,0.00580597794164506,-0.015532210640742,0.00133926835233078,0,-0.028753748665216,-0.0162601287262872,-0.0216064994662132,-0.0115030674846625
"3456",0.00266552297428535,-0.00169287135369067,-0.00390497072230711,-0.00464036007992119,0.00382994042565876,0.000492176633956953,0.00443229283715119,0.00550964168355228,0.00371879985143075,0.00465477114041879
"3457",0.0161669023274218,0.00145350362486374,0.00153402233407429,0.000932360999986281,0,0.00081988263975985,0.0202465640947664,0.00445202039547876,-0.00284997716769297,0
"3458",0.0166093885937895,0.0183841292809257,0.013955137771098,0.0111783572047552,-0.00284643965617914,-0.000163967023723566,0.019972056389937,0.0163654619843165,0.0100605635067958,0.00849420849420857
"3459",-0.00544603705037683,-0.000237520216198384,-0.000839285284608859,-0.000690855578211913,0.0011539615374736,0.000737438722100636,-0.00748317911133922,-0.00939275442444676,0.00843239969041987,-0.0114854517611026
"3460",0.00758201548747262,-0.00546445432371179,-0.00772715502263466,0.0161327454727047,-0.00958515490087586,-0.00270169775895324,0.00326705295314533,0.00609542817150599,-0.00600486552550805,0.0116189000774594
"3461",0.00641991243510498,0.00716672488703574,0.000169343701550417,0.00929912350565476,0.00164957662051801,0.000566797367237637,0.0192886266799359,0.0107708519276624,0.0089205174153264,-0.0122511485451762
"3462",-0.00949437632865391,0.000237182185787388,-0.00490864048884809,-0.0114606435601583,-0.00373419635775518,-0.00098509676560965,0.0159744250383747,0.00133196798761359,-0.000895377743067249,-0.0124031007751938
"3463",0.0177330296912908,0.0175480365178733,0.00816466690333573,0.0134122136845296,-0.0195390567656052,-0.00632754636828048,0.00556362195662019,0.012969704023944,0.00487291942483714,0.0259026687598116
"3464",-0.014215947226743,-0.0144488566814526,-0.0021933958077538,0.00179444972516318,0.00538942602684145,0.00231550180054452,-0.00625441710924479,-0.00755085382635767,-0.011760776729039,0.00382555470543222
"3465",0.0174066610059991,0.00874907384642354,0.00524181154948367,0.0109718543834041,-0.00729288836336306,-0.00288773833025391,0.00108922151504331,0.000661594442606717,-0.000451223906634768,0.00381097560975618
"3466",0.0088625146265493,0.00961089504454771,0.000336454993065338,0.00819483977801649,0.00539992310479276,0.00182050638877196,0.0157176373832881,0.00264462809917343,0.00355493170322241,0.00987091875474566
"3467",0.00893014970480843,0.00928721073921679,-0.000168204677069239,0.00681026241919969,-0.000187365123987315,-0.000495558875390878,-0.00428524229304628,0.00230794592812389,0.0181613488390886,0.00300751879699246
"3468",0.0160876158514391,0.00667125638785593,0.00269090027434937,0.00872786387931734,0.0031857350892539,0.00107423082812397,0.0059773377493535,0.0039473684210527,-0.00287168099324409,-0.0104947526236882
"3469",-0.00652607460337795,-0.0143966877962908,-0.00318682117135016,-0.00410991144142536,0.00716078815584931,0.0022288298076143,-0.01604278273285,-0.0085190039318479,-0.0157288271569432,0.00227272727272743
"3470",-0.00628341482910388,-0.00394162496199124,0.00151433734290518,-0.00673327790077838,0.0022873445558298,0.000329406148885658,-0.0117149999344953,-0.00363516192994062,0.00309477265870606,0.00680272108843538
"3471",-0.001235843736764,-0.0148975484006523,-0.00840052115841949,-0.00721624215883054,-0.00172714913427141,-0.00107034737823641,0.00415488371801631,-0.00132666666666659,0.00364612097052519,0.00300300300300305
"3472",-0.000604308895301053,0.00897925270231559,-0.00203319961696313,0.00352423387864897,-0.00278044039662328,-0.000577014344938287,-0.00620658103418248,-0.0126204246887937,-0.00346520795288618,-0.00673652694610782
"3473",-0.0152034615133015,-0.00538639058369472,0.00118843526105228,-0.00285336324372554,-0.00377967828258707,-0.00164951819869175,-0.0161645934372167,-0.000336394214597968,0.000504744803621726,0.000753579502637436
"3474",0.00400576619007809,0.00824101938340327,0.000169579801137409,0.0110058606741836,-0.00951618289473311,-0.00214781819180598,0.00746827645817838,0.00504717379028174,0.00482090366512078,0.0112951807228916
"3475",-0.00189296396029093,-0.0112096447589269,0.00779921206848044,0.00283048746971337,-0.00345359167253689,-0.00132464494627416,-0.00395353545889299,-0.000334784053070414,0.0075314142259415,-0.00819061801935961
"3476",0.00548533447936417,0.000236078674681561,-0.00285994337268203,-0.000217224939660365,-0.0103968895006082,-0.00348169820447242,-0.00124043760890791,0,-0.00980068627461728,0.00300300300300305
"3477",0.00339515734115792,0.0101535543172981,0.000506113539898934,0.00586323220331564,0.00611254750749457,0.00141420775631906,0.00608552934215889,0.00435361673296653,-0.00106247831949369,-0.00748502994011968
"3478",-0.0184798907440771,-0.0226741371424766,-0.00961217319369589,-0.0129532933979182,0.00930326653020486,0.00265817155273473,-0.0127144919964681,-0.0163387795931976,-0.000503784149707642,-0.0143288084464555
"3479",-0.00344746812040342,-0.0138723282118935,0.00357569448770167,0.00437433195188186,0.00670939990974384,0.00223702136803894,-0.0147536830749667,-0.00813559322033897,0.00263232143434911,0.006885998469778
"3480",-0.0341789145793345,-0.0383215248964798,-0.0135730681597739,-0.0250434789878968,0.000934128924636957,-0.0000826572842642648,-0.0244923785102875,-0.0307586807928913,-0.0161434417128042,-0.026595744680851
"3481",0.0101634726629471,0.00277421491379615,0.00756792706576448,0.0100513889207965,-0.00970741612986192,-0.0042163089676569,0.0152204373609799,0.00846258785392862,-0.0041447282080076,-0.0124902419984387
"3482",-0.0104248295851654,-0.00377261204514623,-0.00580401301547795,-0.011278231774664,-0.00986557732188642,-0.00323787548474364,-0.00679134754081889,-0.00174828671328675,0.00456102068053665,0
"3483",0.0112084430444266,0.0154001473353926,0.0104738204478318,0.0127488167391405,0.00749043717865616,0.00171693127296235,0.0251579592510061,0.00910683044157024,0.00970492071007234,0.0181818181818183
"3484",0.0176559128795439,0.0300844868489389,0.0210705861813798,0.00441692829181006,-0.00580149352506432,-0.00224648270891181,0.0192549505927833,0.0215203409066413,0.00567699385808562,0.0062111801242235
"3485",0.0223491820991495,0.0139994942742572,-0.00166417377804173,0.0314424749755735,0.0216922039246874,0.00842233096993672,0.00209913154406371,0.0142711518858309,-0.000558858714049371,0.0108024691358024
"3486",0.0195028459536541,0.0240420162813715,0.0246708083789295,0.01705391315083,0.00173823997937639,-0.000165380485776523,0.0032034508557035,0.0271356783919598,0.0229839270725449,0.00458015267175571
"3487",-0.00022838487873944,0.00325419373342961,0.000813349375701655,0.00461121750499904,-0.0120847817880022,-0.00339100152029637,-0.00564962190521789,-0.0026092628832356,0.00142135795085285,-0.00379939209726454
"3488",0.0125656639289697,0.029657145342002,0.0294213721099534,0.00688495119009547,-0.0210149548032451,-0.00738586001043107,0.0289031266754562,0.0313931000654022,-0.0442709750065945,0.0122044241037376
"3489",-0.00146660412911126,0.0150765181997541,-0.00378971879777346,-0.0113965383576591,-0.00576692077134833,-0.00284265433565378,0.0111645261366569,0.0174381414889619,0.00331278269005253,0.0195930670685758
"3490",0.00742853389495024,0.00975390288434896,0.00602319847263,0.00649757076191215,0.00360901844252703,0.00159309067793467,0.00641094873379044,0.0137114054222498,-0.00432659673627234,-0.000739098300073904
"3491",-0.00970092595650973,-0.01470905512148,-0.0154403457571992,-0.0074968499512158,0.0170177578901101,0.00569231341892529,-0.0120325176668192,-0.0172148791028243,0.00606068059670717,-0.00813609467455612
"3492",0.013844509855391,0.0155971311749648,0.0142422410626972,0.0140579705290693,-0.00132589186917087,-0.00133172710437202,0.0261492367164731,0.00594310309487334,0.0068197144365878,-0.00447427293064884
"3493",0.0124826120023434,0.00943387302159993,0.0142000283627697,0.0124145558041135,-0.00240269129403659,-0.000750221641979465,0.00814518663445041,0.0130597636815921,-0.0000565025952471432,0.00898876404494398
"3494",-0.00537832385488324,-0.00130399049995145,-0.0038892659950639,-0.0010218603743678,0.00652797809599392,0.00258566754078537,0.000807900658351457,0.00306930613448086,-0.0036691731414904,0.00296956198960641
"3495",-0.0120348718247192,-0.00544065470791644,-0.00671560505874069,-0.003477937055131,0.00289669115395697,-0.000332703138277712,-0.0179909802039316,-0.00489596083231325,-0.0057223512747876,0.00148038490007396
"3496",0.00421022508385915,0.00722093857035078,0.00660374314661683,0.00164244817016623,0.00514840727626309,0.00108191171718053,0.00199648384165196,0.00430504305043033,-0.00188045467318787,0
"3497",-0.00684779803934021,-0.00130342385404636,0.0112465123830972,0.00553387530597993,0.00886997129430211,0.00174571740082841,-0.00468823513752781,-0.00122477036129809,0.00302579349107579,0.00517368810051733
"3498",0.0059943794810573,-0.000870163676983338,0.000617941067318828,0.00264982154223148,-0.00458159322621399,-0.00199168931936677,-0.0008242641758619,-0.00582461697806924,-0.0196938127418315,0.00294117647058822
"3499",0.0161137303668235,0.0156760829074649,0.0151281221610053,0.013417310619622,-0.00995223795148559,-0.00157990938871044,0.00282848676865965,0.0141843663274748,-0.015328340366448,0.0212609970674487
"3500",-0.00154174863315815,0.000214267322909523,-0.00714722697049641,-0.00561683332116936,-0.00307851511692148,0.000333121714970908,0.000822712080600807,0.00121620557057467,-0.000471731834936873,0.00861450107681261
"3501",0.00278504414703007,0.00364340506008598,0.014397339729274,0.00948162992926993,0.00970510441013284,0.00299726376293741,-0.00305307807835509,0.00182210750075917,-0.0101469060865702,-0.0021352313167261
"3502",-0.00442712815826585,-0.0164424191356956,-0.0277819728086511,-0.0261790905105282,-0.00124816437080588,-0.000664039598186839,-0.00871616470103909,-0.017278083220486,-0.00667498090902252,-0.00570613409415122
"3503",0.0109373702926832,0.0245331782243872,0.020500059348493,0.0197003132712501,-0.0147444903241852,-0.00531958933512211,0.0114069099515917,0.021283252392551,0.0210595490617334,-0.00286944045911042
"3504",0.00210377143133078,0.0012714691306086,-0.00167407295458155,0.00140878066887606,-0.007936543347558,-0.00167123596585095,-0.00892862287981588,-0.00634246432067442,0.00752153045393533,0.00431654676258986
"3505",-0.00027264501842017,0.000846591020783549,0.00243908452286878,0.0114550570768115,0.00806397460988029,0.00267846224921109,0.00746790859911606,0.0103343458763314,0.00787350370281992,0.00143266475644688
"3506",0.00861760247602539,0.00888127115526061,0.00456194608143701,0.0103317284283577,-0.014665699235193,-0.00392350993706891,0.0147076629402403,0.00661844123836119,-0.0028354320101317,0.0042918454935621
"3507",-0.00205488945832433,-0.00523993063764894,-0.0146835712894194,0,0.00902063734986602,0.0031008996176265,-0.00776899176447665,-0.00717268401591997,0.014914066246527,0
"3508",0.0029261812179262,0.00400338131424816,0.00230451390225084,0.000393286902139467,0.00472540948529798,0.00100258237316964,-0.00490830012383747,0.00361225154689193,0.00348791242202484,0.00142450142450157
"3509",-0.00896893548350419,-0.000419689281515145,0.00705086648059527,-0.00864948631826545,-0.00330492482629707,-0.00141893447666108,-0.00763353884671281,-0.0026994601079785,-0.0170940170940171,0.000711237553342903
"3510",-0.000327069065734764,-0.00125980799217373,0.00167422087668445,0.0128892379962506,0.00886364905207349,0.00225684097078482,-0.00579881358040146,0.00330830075187971,-0.00191305507246387,0.0149253731343284
"3511",-0.00117257171203444,-0.0060962691463915,0.00212740790044719,-0.00704776281654174,0.00353960911229589,0.00200149411314832,0.000476098068984854,0.000599520365721862,0.00185866877921437,-0.00280112044817926
"3512",-0.00447716915727869,-0.000681773644459427,0.00331856233150818,-0.00519919880486852,-0.00277132019028492,-0.000582643638787683,-0.00466151798085734,0.00149787293295756,-0.0055076350655795,0.00280898876404478
"3513",0.0135193949138301,0.0138592104964088,0.00713082948682575,0.0108129958112333,-0.0033474534180945,-0.000999326155221913,0.0192632559418073,0.010768800478612,0.0139909589479812,0.00770308123249319
"3514",0.0015694094177825,0.00462672985545187,-0.000150557403610696,0.00475437797147404,-0.00266155683820046,-0.000833593717547543,0.00153551847221745,0.00680671776245312,0.00551909847626653,0.00555941626129264
"3515",0.00559195502136389,0.00795482520410284,0.00587613352978167,0.00650626958780998,-0.00264604106491628,-0.00072633923398191,0.0097889136715541,0.00646684303350953,0.0105203605667363,0.0117484450587422
"3516",-0.00399290720344347,-0.00373833837016246,-0.00284604545098732,-0.0011752595724831,-0.00299745529979356,-0.000835413554772235,-0.0179864628129014,-0.0140188075923592,-0.00169742554890162,0.00341530054644812
